
module SK_gen_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module SK_gen_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module SK_gen_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  TIE0DHD U1 ( .O(n1) );
endmodule


module SK_gen_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_add_8 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_add_6 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_add_5 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  INVDHD U1 ( .I(B[4]), .O(n4) );
  INVDHD U2 ( .I(B[3]), .O(n5) );
  INVDHD U3 ( .I(B[2]), .O(n6) );
  INVDHD U4 ( .I(B[5]), .O(n3) );
  INVDHD U5 ( .I(B[6]), .O(n2) );
  INVDHD U6 ( .I(B[1]), .O(n7) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_add_4 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_sub_6 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  INVDHD U1 ( .I(B[3]), .O(n5) );
  INVDHD U2 ( .I(B[2]), .O(n6) );
  INVDHD U3 ( .I(B[4]), .O(n4) );
  INVDHD U4 ( .I(B[5]), .O(n3) );
  INVDHD U5 ( .I(B[6]), .O(n2) );
  INVDHD U6 ( .I(B[1]), .O(n7) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVDHD U1 ( .I(B[2]), .O(n6) );
  INVDHD U2 ( .I(B[5]), .O(n3) );
  INVDHD U3 ( .I(B[1]), .O(n7) );
  INVDHD U4 ( .I(B[3]), .O(n5) );
  INVDHD U5 ( .I(B[4]), .O(n4) );
  INVDHD U6 ( .I(B[6]), .O(n2) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_sub_4 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVDHD U1 ( .I(B[2]), .O(n6) );
  INVDHD U2 ( .I(B[3]), .O(n5) );
  INVDHD U3 ( .I(B[4]), .O(n4) );
  INVDHD U4 ( .I(B[5]), .O(n3) );
  INVDHD U5 ( .I(B[6]), .O(n2) );
  INVDHD U6 ( .I(B[1]), .O(n7) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_sub_3 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVDHD U1 ( .I(B[2]), .O(n6) );
  INVDHD U2 ( .I(B[5]), .O(n3) );
  INVDHD U3 ( .I(B[1]), .O(n7) );
  INVDHD U4 ( .I(B[3]), .O(n5) );
  INVDHD U5 ( .I(B[4]), .O(n4) );
  INVDHD U6 ( .I(B[6]), .O(n2) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_sub_2 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVDHD U1 ( .I(B[2]), .O(n6) );
  INVDHD U2 ( .I(B[5]), .O(n3) );
  INVDHD U3 ( .I(B[1]), .O(n7) );
  INVDHD U4 ( .I(B[3]), .O(n5) );
  INVDHD U5 ( .I(B[4]), .O(n4) );
  INVDHD U6 ( .I(B[6]), .O(n2) );
  INVDHD U7 ( .I(B[0]), .O(n8) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  INVDHD U1 ( .I(B[7]), .O(n1) );
  INVDHD U2 ( .I(B[5]), .O(n3) );
  INVDHD U3 ( .I(B[3]), .O(n5) );
  INVDHD U4 ( .I(B[4]), .O(n4) );
  INVDHD U5 ( .I(B[6]), .O(n2) );
  INVDHD U6 ( .I(B[1]), .O(n7) );
  INVDHD U7 ( .I(B[2]), .O(n6) );
  INVDHD U8 ( .I(B[0]), .O(n8) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [8:0] carry;

  FA1DHD U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FA1DHD U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FA1DHD U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FA1DHD U2_0 ( .A(A[0]), .B(n8), .CI(n9), .CO(carry[1]), .S(DIFF[0]) );
  FA1DHD U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FA1DHD U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FA1DHD U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  XOR3EHD U2_7 ( .I1(A[7]), .I2(n1), .I3(carry[7]), .O(DIFF[7]) );
  INVDHD U1 ( .I(B[2]), .O(n6) );
  INVDHD U2 ( .I(B[1]), .O(n7) );
  INVDHD U3 ( .I(B[5]), .O(n3) );
  INVDHD U4 ( .I(B[0]), .O(n8) );
  INVDHD U5 ( .I(B[3]), .O(n5) );
  INVDHD U6 ( .I(B[4]), .O(n4) );
  INVDHD U7 ( .I(B[6]), .O(n2) );
  INVDHD U8 ( .I(B[7]), .O(n1) );
  TIE1DHD U9 ( .O(n9) );
endmodule


module round_funct_DW01_add_0 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [7:1] carry;

  XOR3EHD U1_7 ( .I1(A[7]), .I2(B[7]), .I3(carry[7]), .O(SUM[7]) );
  FA1DHD U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FA1DHD U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FA1DHD U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FA1DHD U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FA1DHD U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FA1DHD U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(SUM[1])
         );
  FA1DHD U1_0 ( .A(A[0]), .B(B[0]), .CI(n1), .CO(carry[1]), .S(SUM[0]) );
  TIE0DHD U1 ( .O(n1) );
endmodule


module round_funct ( P, MK, SKx0, SKx1, SKx2, SKx3, clk, reset, ed, WK0_4, 
        WK1_5, WK2_6, WK3_7, C );
  input [63:0] P;
  input [127:0] MK;
  input [7:0] SKx0;
  input [7:0] SKx1;
  input [7:0] SKx2;
  input [7:0] SKx3;
  input [7:0] WK0_4;
  input [7:0] WK1_5;
  input [7:0] WK2_6;
  input [7:0] WK3_7;
  output [63:0] C;
  input clk, reset, ed;
  wire   N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N23, N26, N27, N28, N29, N30, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N75, N76, N77, N78, N79,
         N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N173, N174, N175,
         N176, N177, N178, N179, N180, N197, N198, N199, N200, N201, N202,
         N203, N204, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, N266, N267, N268, N269, N270, N287, N288, N289, N290,
         N291, N292, N293, N294, N295, N296, N297, N298, N299, N300, N301,
         N302, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N412, N421, N422, N423, N424, N425, N426, N427, N428,
         N429, N430, N431, N432, N433, N434, N435, N436, N437, N438, N439,
         N440, N441, N442, N443, N444, n1, n171, n172, n173, n174, n175, n176,
         n177, n178, n182, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, \add_49/carry[5] ,
         \add_49/carry[4] , \add_49/carry[3] , \add_49/carry[2] , n2, n3, n4,
         n5, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n179, n180, n181, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332;
  wire   [7:0] X6x;
  wire   [7:0] X2x;
  wire   [7:0] X3x;
  wire   [7:0] X7x;
  wire   [7:0] X0x;
  wire   [7:0] X4x;
  wire   [7:0] X5x;
  wire   [7:0] X1x;
  wire   [7:0] F0X6;
  wire   [7:0] F0X2;
  wire   [7:0] F0X3;
  wire   [7:0] F0X7;
  wire   [5:0] i_round;
  wire   [7:0] X00x;

  round_funct_DW01_add_0 add_121 ( .A(F0X7), .B(SKx3), .CI(n1), .SUM({N444, 
        N443, N442, N441, N440, N439, N438, N437}) );
  round_funct_DW01_sub_0 sub_119 ( .A(X6x), .B({N421, N422, N423, N424, N425, 
        N426, N427, N428}), .CI(n1), .DIFF({N436, N435, N434, N433, N432, N431, 
        N430, N429}) );
  round_funct_DW01_add_1 add_117 ( .A(F0X3), .B(SKx1), .CI(n1), .SUM({N412, 
        N411, N410, N409, N408, N407, N406, N405}) );
  round_funct_DW01_sub_1 sub_115 ( .A(X2x), .B({N389, N390, N391, N392, N393, 
        N394, N395, N396}), .CI(n1), .DIFF({N404, N403, N402, N401, N400, N399, 
        N398, N397}) );
  round_funct_DW01_sub_2 sub_106 ( .A(X4x), .B(WK2_6), .CI(n1), .DIFF({N302, 
        N301, N300, N299, N298, N297, N296, N295}) );
  round_funct_DW01_add_2 add_106 ( .A(X4x), .B(WK2_6), .CI(n1), .SUM({N294, 
        N293, N292, N291, N290, N289, N288, N287}) );
  round_funct_DW01_sub_3 sub_102 ( .A(X0x), .B(WK0_4), .CI(n1), .DIFF({N270, 
        N269, N268, N267, N266, N265, N264, N263}) );
  round_funct_DW01_add_3 add_102 ( .A(X0x), .B(WK0_4), .CI(n1), .SUM({N262, 
        N261, N260, N259, N258, N257, N256, N255}) );
  round_funct_DW01_sub_4 sub_70 ( .A(X5x), .B({N14, N15, N16, N17, N18, N19, 
        N20, N21}), .CI(n1), .DIFF({N139, N138, N137, N136, N135, N134, N133, 
        N132}) );
  round_funct_DW01_sub_5 sub_66 ( .A(X1x), .B({N6, N7, N8, N9, N10, N11, N12, 
        N13}), .CI(n1), .DIFF({N115, N114, N113, N112, N111, N110, N109, N108}) );
  round_funct_DW01_sub_6 sub_57 ( .A(P[39:32]), .B(WK2_6), .CI(n1), .DIFF({N90, 
        N89, N88, N87, N86, N85, N84, N83}) );
  round_funct_DW01_add_4 add_57 ( .A(P[39:32]), .B(WK2_6), .CI(n1), .SUM({N82, 
        N81, N80, N79, N78, N77, N76, N75}) );
  round_funct_DW01_sub_7 sub_53 ( .A(P[7:0]), .B(WK0_4), .CI(n1), .DIFF({N58, 
        N57, N56, N55, N54, N53, N52, N51}) );
  round_funct_DW01_add_5 add_53 ( .A(P[7:0]), .B(WK0_4), .CI(n1), .SUM({N50, 
        N49, N48, N47, N46, N45, N44, N43}) );
  round_funct_DW01_add_6 r138 ( .A(X5x), .B({N14, N15, N16, N17, N18, N19, N20, 
        N21}), .CI(n1), .SUM({N204, N203, N202, N201, N200, N199, N198, N197})
         );
  round_funct_DW01_add_7 r137 ( .A(X1x), .B({N6, N7, N8, N9, N10, N11, N12, 
        N13}), .CI(n1), .SUM({N180, N179, N178, N177, N176, N175, N174, N173})
         );
  round_funct_DW01_add_8 r136 ( .A(F0X6), .B(SKx3), .CI(n1), .SUM({N147, N146, 
        N145, N144, N143, N142, N141, N140}) );
  round_funct_DW01_add_9 r134 ( .A(F0X2), .B(SKx1), .CI(n1), .SUM({N123, N122, 
        N121, N120, N119, N118, N117, N116}) );
  DFECHD \X00x_reg[7]  ( .D(X0x[7]), .EB(n315), .CK(clk), .Q(X00x[7]) );
  DFECHD \X00x_reg[0]  ( .D(X0x[0]), .EB(n315), .CK(clk), .Q(X00x[0]) );
  DFECHD \X00x_reg[1]  ( .D(X0x[1]), .EB(n315), .CK(clk), .Q(X00x[1]) );
  DFECHD \X00x_reg[2]  ( .D(X0x[2]), .EB(n315), .CK(clk), .Q(X00x[2]) );
  DFECHD \X00x_reg[3]  ( .D(X0x[3]), .EB(n315), .CK(clk), .Q(X00x[3]) );
  DFECHD \X00x_reg[4]  ( .D(X0x[4]), .EB(n315), .CK(clk), .Q(X00x[4]) );
  DFECHD \X00x_reg[5]  ( .D(X0x[5]), .EB(n315), .CK(clk), .Q(X00x[5]) );
  DFECHD \X00x_reg[6]  ( .D(X0x[6]), .EB(n315), .CK(clk), .Q(X00x[6]) );
  QDFFEHD \C0_reg[0]  ( .D(n407), .CK(clk), .Q(C[0]) );
  QDFFEHD \C0_reg[1]  ( .D(n406), .CK(clk), .Q(C[1]) );
  QDFFEHD \C0_reg[2]  ( .D(n405), .CK(clk), .Q(C[2]) );
  QDFFEHD \C0_reg[3]  ( .D(n404), .CK(clk), .Q(C[3]) );
  QDFFEHD \C0_reg[4]  ( .D(n403), .CK(clk), .Q(C[4]) );
  QDFFEHD \C0_reg[5]  ( .D(n402), .CK(clk), .Q(C[5]) );
  QDFFEHD \C0_reg[6]  ( .D(n401), .CK(clk), .Q(C[6]) );
  QDFFEHD \C0_reg[7]  ( .D(n400), .CK(clk), .Q(C[7]) );
  QDFFEHD \C4_reg[7]  ( .D(n375), .CK(clk), .Q(C[39]) );
  QDFFEHD \C4_reg[6]  ( .D(n374), .CK(clk), .Q(C[38]) );
  QDFFEHD \C4_reg[5]  ( .D(n373), .CK(clk), .Q(C[37]) );
  QDFFEHD \C4_reg[4]  ( .D(n372), .CK(clk), .Q(C[36]) );
  QDFFEHD \C4_reg[3]  ( .D(n371), .CK(clk), .Q(C[35]) );
  QDFFEHD \C4_reg[2]  ( .D(n370), .CK(clk), .Q(C[34]) );
  QDFFEHD \C4_reg[1]  ( .D(n369), .CK(clk), .Q(C[33]) );
  QDFFEHD \C4_reg[0]  ( .D(n368), .CK(clk), .Q(C[32]) );
  DFCLRBEHD \i_round_reg[0]  ( .RB(n332), .D(n5), .LD(N23), .CK(clk), .Q(n306), 
        .QB(n5) );
  QDFFEHD \X3x_reg[6]  ( .D(n377), .CK(clk), .Q(X3x[6]) );
  QDFFEHD \X3x_reg[5]  ( .D(n378), .CK(clk), .Q(X3x[5]) );
  QDFFEHD \X3x_reg[1]  ( .D(n382), .CK(clk), .Q(X3x[1]) );
  QDFFEHD \X3x_reg[2]  ( .D(n381), .CK(clk), .Q(X3x[2]) );
  QDFFEHD \X3x_reg[3]  ( .D(n380), .CK(clk), .Q(X3x[3]) );
  QDFFEHD \X3x_reg[4]  ( .D(n379), .CK(clk), .Q(X3x[4]) );
  QDFFEHD \X3x_reg[0]  ( .D(n383), .CK(clk), .Q(X3x[0]) );
  QDFFEHD \X7x_reg[3]  ( .D(n420), .CK(clk), .Q(X7x[3]) );
  QDFFEHD \X7x_reg[4]  ( .D(n419), .CK(clk), .Q(X7x[4]) );
  QDFFEHD \X7x_reg[0]  ( .D(n423), .CK(clk), .Q(X7x[0]) );
  QDFFEHD \X7x_reg[5]  ( .D(n418), .CK(clk), .Q(X7x[5]) );
  QDFFEHD \X7x_reg[2]  ( .D(n421), .CK(clk), .Q(X7x[2]) );
  QDFFEHD \X6x_reg[4]  ( .D(n427), .CK(clk), .Q(X6x[4]) );
  QDFFEHD \X6x_reg[5]  ( .D(n426), .CK(clk), .Q(X6x[5]) );
  QDFFEHD \X4x_reg[7]  ( .D(n439), .CK(clk), .Q(X4x[7]) );
  QDFFEHD \X4x_reg[0]  ( .D(n446), .CK(clk), .Q(X4x[0]) );
  QDFFEHD \X1x_reg[7]  ( .D(n392), .CK(clk), .Q(X1x[7]) );
  QDFFEHD \X1x_reg[0]  ( .D(n399), .CK(clk), .Q(X1x[0]) );
  QDFFEHD \X0x_reg[7]  ( .D(n408), .CK(clk), .Q(X0x[7]) );
  QDFFEHD \X0x_reg[0]  ( .D(n415), .CK(clk), .Q(X0x[0]) );
  QDFFEHD \X2x_reg[4]  ( .D(n387), .CK(clk), .Q(X2x[4]) );
  QDFFEHD \X4x_reg[1]  ( .D(n445), .CK(clk), .Q(X4x[1]) );
  QDFFEHD \X1x_reg[6]  ( .D(n393), .CK(clk), .Q(X1x[6]) );
  QDFFEHD \X1x_reg[3]  ( .D(n396), .CK(clk), .Q(X1x[3]) );
  QDFFEHD \X1x_reg[4]  ( .D(n395), .CK(clk), .Q(X1x[4]) );
  QDFFEHD \X1x_reg[1]  ( .D(n398), .CK(clk), .Q(X1x[1]) );
  QDFFEHD \X0x_reg[1]  ( .D(n414), .CK(clk), .Q(X0x[1]) );
  QDFFEHD \X2x_reg[5]  ( .D(n386), .CK(clk), .Q(X2x[5]) );
  QDFFEHD \X3x_reg[7]  ( .D(n376), .CK(clk), .Q(X3x[7]) );
  QDFFEHD \X7x_reg[7]  ( .D(n416), .CK(clk), .Q(X7x[7]) );
  QDFFEHD \X7x_reg[6]  ( .D(n417), .CK(clk), .Q(X7x[6]) );
  QDFFEHD \X6x_reg[7]  ( .D(n424), .CK(clk), .Q(X6x[7]) );
  QDFFEHD \X7x_reg[1]  ( .D(n422), .CK(clk), .Q(X7x[1]) );
  QDFFEHD \X6x_reg[6]  ( .D(n425), .CK(clk), .Q(X6x[6]) );
  QDFFEHD \X2x_reg[0]  ( .D(n391), .CK(clk), .Q(X2x[0]) );
  QDFFEHD \X2x_reg[1]  ( .D(n390), .CK(clk), .Q(X2x[1]) );
  QDFFEHD \X2x_reg[2]  ( .D(n389), .CK(clk), .Q(X2x[2]) );
  QDFFEHD \X6x_reg[3]  ( .D(n428), .CK(clk), .Q(X6x[3]) );
  QDFFEHD \X6x_reg[0]  ( .D(n431), .CK(clk), .Q(X6x[0]) );
  QDFFEHD \X6x_reg[1]  ( .D(n430), .CK(clk), .Q(X6x[1]) );
  QDFFEHD \X6x_reg[2]  ( .D(n429), .CK(clk), .Q(X6x[2]) );
  QDFFEHD \X2x_reg[7]  ( .D(n384), .CK(clk), .Q(X2x[7]) );
  QDFFEHD \X2x_reg[6]  ( .D(n385), .CK(clk), .Q(X2x[6]) );
  QDFFEHD \X2x_reg[3]  ( .D(n388), .CK(clk), .Q(X2x[3]) );
  QDFFEHD \X4x_reg[6]  ( .D(n440), .CK(clk), .Q(X4x[6]) );
  QDFFEHD \X4x_reg[4]  ( .D(n442), .CK(clk), .Q(X4x[4]) );
  QDFFEHD \X4x_reg[3]  ( .D(n443), .CK(clk), .Q(X4x[3]) );
  QDFFEHD \X0x_reg[6]  ( .D(n409), .CK(clk), .Q(X0x[6]) );
  QDFFEHD \X0x_reg[3]  ( .D(n412), .CK(clk), .Q(X0x[3]) );
  QDFFEHD \X0x_reg[4]  ( .D(n411), .CK(clk), .Q(X0x[4]) );
  QDFFEHD \X4x_reg[5]  ( .D(n441), .CK(clk), .Q(X4x[5]) );
  QDFFEHD \X4x_reg[2]  ( .D(n444), .CK(clk), .Q(X4x[2]) );
  QDFFEHD \X1x_reg[5]  ( .D(n394), .CK(clk), .Q(X1x[5]) );
  QDFFEHD \X1x_reg[2]  ( .D(n397), .CK(clk), .Q(X1x[2]) );
  QDFFEHD \X0x_reg[5]  ( .D(n410), .CK(clk), .Q(X0x[5]) );
  QDFFEHD \X0x_reg[2]  ( .D(n413), .CK(clk), .Q(X0x[2]) );
  DFECHD \C2_reg[7]  ( .D(n316), .EB(n102), .CK(clk), .Q(C[23]) );
  DFECHD \C6_reg[6]  ( .D(n318), .EB(n101), .CK(clk), .Q(C[54]) );
  DFECHD \C2_reg[0]  ( .D(n319), .EB(n101), .CK(clk), .Q(C[16]) );
  DFECHD \C6_reg[0]  ( .D(n321), .EB(n101), .CK(clk), .Q(C[48]) );
  DFECHD \C6_reg[1]  ( .D(n322), .EB(n101), .CK(clk), .Q(C[49]) );
  DFECHD \C2_reg[1]  ( .D(n323), .EB(n100), .CK(clk), .Q(C[17]) );
  DFECHD \C6_reg[2]  ( .D(n324), .EB(n100), .CK(clk), .Q(C[50]) );
  DFECHD \C2_reg[2]  ( .D(n325), .EB(n100), .CK(clk), .Q(C[18]) );
  DFECHD \C6_reg[3]  ( .D(n326), .EB(n99), .CK(clk), .Q(C[51]) );
  DFECHD \C2_reg[3]  ( .D(n327), .EB(n99), .CK(clk), .Q(C[19]) );
  DFECHD \C6_reg[4]  ( .D(n328), .EB(n99), .CK(clk), .Q(C[52]) );
  DFECHD \C6_reg[7]  ( .D(n329), .EB(n99), .CK(clk), .Q(C[55]) );
  DFECHD \C2_reg[4]  ( .D(n330), .EB(n99), .CK(clk), .Q(C[20]) );
  DFECHD \C2_reg[5]  ( .D(n320), .EB(n98), .CK(clk), .Q(C[21]) );
  DFECHD \C6_reg[5]  ( .D(n331), .EB(n98), .CK(clk), .Q(C[53]) );
  DFECHD \C2_reg[6]  ( .D(n317), .EB(n98), .CK(clk), .Q(C[22]) );
  DFECHD \C3_reg[0]  ( .D(X3x[0]), .EB(n102), .CK(clk), .Q(C[24]) );
  DFECHD \C3_reg[7]  ( .D(X3x[7]), .EB(n102), .CK(clk), .Q(C[31]) );
  DFECHD \C3_reg[6]  ( .D(X3x[6]), .EB(n102), .CK(clk), .Q(C[30]) );
  DFECHD \C7_reg[7]  ( .D(X7x[7]), .EB(n101), .CK(clk), .Q(C[63]) );
  DFECHD \C7_reg[6]  ( .D(X7x[6]), .EB(n101), .CK(clk), .Q(C[62]) );
  DFECHD \C7_reg[0]  ( .D(X7x[0]), .EB(n101), .CK(clk), .Q(C[56]) );
  DFECHD \C1_reg[0]  ( .D(X1x[0]), .EB(n101), .CK(clk), .Q(C[8]) );
  DFECHD \C7_reg[1]  ( .D(X7x[1]), .EB(n101), .CK(clk), .Q(C[57]) );
  DFECHD \C1_reg[1]  ( .D(X1x[1]), .EB(n101), .CK(clk), .Q(C[9]) );
  DFECHD \C3_reg[1]  ( .D(X3x[1]), .EB(n100), .CK(clk), .Q(C[25]) );
  DFECHD \C5_reg[1]  ( .D(X5x[1]), .EB(n100), .CK(clk), .Q(C[41]) );
  DFECHD \C7_reg[2]  ( .D(X7x[2]), .EB(n100), .CK(clk), .Q(C[58]) );
  DFECHD \C1_reg[2]  ( .D(X1x[2]), .EB(n100), .CK(clk), .Q(C[10]) );
  DFECHD \C3_reg[2]  ( .D(X3x[2]), .EB(n100), .CK(clk), .Q(C[26]) );
  DFECHD \C5_reg[2]  ( .D(X5x[2]), .EB(n100), .CK(clk), .Q(C[42]) );
  DFECHD \C7_reg[3]  ( .D(X7x[3]), .EB(n100), .CK(clk), .Q(C[59]) );
  DFECHD \C1_reg[3]  ( .D(X1x[3]), .EB(n100), .CK(clk), .Q(C[11]) );
  DFECHD \C3_reg[3]  ( .D(X3x[3]), .EB(n99), .CK(clk), .Q(C[27]) );
  DFECHD \C5_reg[3]  ( .D(X5x[3]), .EB(n99), .CK(clk), .Q(C[43]) );
  DFECHD \C7_reg[4]  ( .D(X7x[4]), .EB(n99), .CK(clk), .Q(C[60]) );
  DFECHD \C1_reg[4]  ( .D(X1x[4]), .EB(n99), .CK(clk), .Q(C[12]) );
  DFECHD \C3_reg[4]  ( .D(X3x[4]), .EB(n99), .CK(clk), .Q(C[28]) );
  DFECHD \C5_reg[4]  ( .D(X5x[4]), .EB(n99), .CK(clk), .Q(C[44]) );
  DFECHD \C5_reg[5]  ( .D(X5x[5]), .EB(n98), .CK(clk), .Q(C[45]) );
  DFECHD \C3_reg[5]  ( .D(X3x[5]), .EB(n98), .CK(clk), .Q(C[29]) );
  DFECHD \C7_reg[5]  ( .D(X7x[5]), .EB(n98), .CK(clk), .Q(C[61]) );
  DFECHD \C1_reg[5]  ( .D(X1x[5]), .EB(n98), .CK(clk), .Q(C[13]) );
  DFECHD \C1_reg[6]  ( .D(X1x[6]), .EB(n98), .CK(clk), .Q(C[14]) );
  DFECHD \C1_reg[7]  ( .D(X1x[7]), .EB(n98), .CK(clk), .Q(C[15]) );
  DFECHD \C5_reg[6]  ( .D(X5x[6]), .EB(n98), .CK(clk), .Q(C[46]) );
  DFECHD \C5_reg[7]  ( .D(X5x[7]), .EB(n98), .CK(clk), .Q(C[47]) );
  DFECHD \C5_reg[0]  ( .D(X5x[0]), .EB(n101), .CK(clk), .Q(C[40]) );
  DFCLRBEHD \i_round_reg[5]  ( .RB(n332), .D(N30), .LD(N23), .CK(clk), .Q(
        i_round[5]), .QB(n108) );
  DFCLRBEHD \i_round_reg[4]  ( .RB(n332), .D(N29), .LD(N23), .CK(clk), .Q(
        i_round[4]), .QB(n104) );
  DFCLRBEHD \i_round_reg[3]  ( .RB(n332), .D(N28), .LD(N23), .CK(clk), .Q(
        i_round[3]), .QB(n105) );
  DFCLRBEHD \i_round_reg[2]  ( .RB(n332), .D(N27), .LD(N23), .CK(clk), .Q(
        i_round[2]), .QB(n106) );
  DFCLRBEHD \i_round_reg[1]  ( .RB(n332), .D(N26), .LD(N23), .CK(clk), .Q(n311), .QB(n107) );
  DFFCHD \X5x_reg[7]  ( .D(n432), .CK(clk), .Q(X5x[7]), .QB(n171) );
  DFFCHD \X5x_reg[4]  ( .D(n435), .CK(clk), .Q(X5x[4]), .QB(n174) );
  DFFCHD \X5x_reg[3]  ( .D(n436), .CK(clk), .Q(X5x[3]), .QB(n175) );
  DFFCHD \X5x_reg[6]  ( .D(n433), .CK(clk), .Q(X5x[6]), .QB(n172) );
  DFFCHD \X5x_reg[5]  ( .D(n434), .CK(clk), .Q(X5x[5]), .QB(n173) );
  DFFCHD \X5x_reg[1]  ( .D(n438), .CK(clk), .Q(X5x[1]), .QB(n177) );
  DFFCHD \X5x_reg[0]  ( .D(n447), .CK(clk), .Q(X5x[0]), .QB(n178) );
  DFFCHD \X5x_reg[2]  ( .D(n437), .CK(clk), .Q(X5x[2]), .QB(n176) );
  AN3EHD U3 ( .I1(n108), .I2(n246), .I3(n305), .O(n2) );
  OA112EHD U4 ( .C1(n306), .C2(n308), .A1(n246), .B1(n309), .O(n3) );
  AN2EHD U5 ( .I1(ed), .I2(n309), .O(n4) );
  INVDHD U6 ( .I(n63), .O(n113) );
  INVDHD U7 ( .I(n62), .O(n179) );
  BUFEHD U8 ( .I(n112), .O(n62) );
  NR2CHD U9 ( .I1(n113), .I2(n76), .O(n112) );
  BUFEHD U10 ( .I(n162), .O(n63) );
  NR3BHD U11 ( .I1(n90), .I2(n71), .I3(n82), .O(n162) );
  BUFEHD U12 ( .I(n96), .O(n103) );
  BUFEHD U13 ( .I(n78), .O(n80) );
  BUFEHD U14 ( .I(n78), .O(n81) );
  BUFEHD U15 ( .I(n78), .O(n82) );
  BUFEHD U16 ( .I(n79), .O(n83) );
  BUFEHD U17 ( .I(n79), .O(n84) );
  BUFEHD U18 ( .I(n94), .O(n98) );
  BUFEHD U19 ( .I(n94), .O(n99) );
  BUFEHD U20 ( .I(n95), .O(n100) );
  BUFEHD U21 ( .I(n95), .O(n101) );
  BUFEHD U22 ( .I(n96), .O(n102) );
  BUFEHD U23 ( .I(n66), .O(n71) );
  BUFEHD U24 ( .I(n111), .O(n78) );
  BUFEHD U25 ( .I(n2), .O(n76) );
  BUFEHD U26 ( .I(n97), .O(n96) );
  BUFEHD U27 ( .I(n77), .O(n74) );
  BUFEHD U28 ( .I(n77), .O(n75) );
  BUFEHD U29 ( .I(n85), .O(n88) );
  BUFEHD U30 ( .I(n65), .O(n68) );
  BUFEHD U31 ( .I(n85), .O(n89) );
  BUFEHD U32 ( .I(n65), .O(n69) );
  BUFEHD U33 ( .I(n86), .O(n90) );
  BUFEHD U34 ( .I(n66), .O(n70) );
  BUFEHD U35 ( .I(n86), .O(n91) );
  BUFEHD U36 ( .I(n87), .O(n92) );
  BUFEHD U37 ( .I(n67), .O(n72) );
  BUFEHD U38 ( .I(n67), .O(n73) );
  BUFEHD U39 ( .I(n111), .O(n79) );
  BUFEHD U40 ( .I(n87), .O(n93) );
  BUFEHD U41 ( .I(n97), .O(n94) );
  BUFEHD U42 ( .I(n97), .O(n95) );
  BUFEHD U43 ( .I(n3), .O(n66) );
  NR2CHD U44 ( .I1(n246), .I2(n103), .O(n247) );
  NR2CHD U45 ( .I1(n245), .I2(n246), .O(n119) );
  BUFEHD U46 ( .I(n182), .O(n97) );
  BUFEHD U47 ( .I(n3), .O(n65) );
  BUFEHD U48 ( .I(n3), .O(n67) );
  BUFEHD U49 ( .I(n4), .O(n86) );
  BUFEHD U50 ( .I(n4), .O(n85) );
  BUFEHD U51 ( .I(n4), .O(n87) );
  BUFEHD U52 ( .I(n2), .O(n77) );
  NR2CHD U53 ( .I1(n245), .I2(ed), .O(n117) );
  BUFEHD U54 ( .I(n248), .O(n64) );
  NR2CHD U55 ( .I1(n103), .I2(ed), .O(n248) );
  HA1EHD U56 ( .A(n311), .B(n306), .C(\add_49/carry[2] ), .S(N26) );
  HA1EHD U57 ( .A(i_round[2]), .B(\add_49/carry[2] ), .C(\add_49/carry[3] ), 
        .S(N27) );
  HA1EHD U58 ( .A(i_round[3]), .B(\add_49/carry[3] ), .C(\add_49/carry[4] ), 
        .S(N28) );
  HA1EHD U59 ( .A(i_round[4]), .B(\add_49/carry[4] ), .C(\add_49/carry[5] ), 
        .S(N29) );
  TIE0DHD U60 ( .O(n1) );
  XOR2CHD U61 ( .I1(\add_49/carry[5] ), .I2(i_round[5]), .O(N30) );
  NR2BHD U62 ( .I1(n71), .I2(n77), .O(n315) );
  XOR2CHD U63 ( .I1(X2x[7]), .I2(WK1_5[7]), .O(n316) );
  XOR2CHD U64 ( .I1(X2x[6]), .I2(WK1_5[6]), .O(n317) );
  XOR2CHD U65 ( .I1(X6x[6]), .I2(WK3_7[6]), .O(n318) );
  XOR2CHD U66 ( .I1(X2x[0]), .I2(WK1_5[0]), .O(n319) );
  XOR2CHD U67 ( .I1(X2x[5]), .I2(WK1_5[5]), .O(n320) );
  XOR2CHD U68 ( .I1(X6x[0]), .I2(WK3_7[0]), .O(n321) );
  XOR2CHD U69 ( .I1(X6x[1]), .I2(WK3_7[1]), .O(n322) );
  XOR2CHD U70 ( .I1(X2x[1]), .I2(WK1_5[1]), .O(n323) );
  XOR2CHD U71 ( .I1(X6x[2]), .I2(WK3_7[2]), .O(n324) );
  XOR2CHD U72 ( .I1(X2x[2]), .I2(WK1_5[2]), .O(n325) );
  XOR2CHD U73 ( .I1(X6x[3]), .I2(WK3_7[3]), .O(n326) );
  XOR2CHD U74 ( .I1(X2x[3]), .I2(WK1_5[3]), .O(n327) );
  XOR2CHD U75 ( .I1(X6x[4]), .I2(WK3_7[4]), .O(n328) );
  XOR2CHD U76 ( .I1(X6x[7]), .I2(WK3_7[7]), .O(n329) );
  XOR2CHD U77 ( .I1(X2x[4]), .I2(WK1_5[4]), .O(n330) );
  XOR2CHD U78 ( .I1(X6x[5]), .I2(WK3_7[5]), .O(n331) );
  INVCHD U79 ( .I(reset), .O(n332) );
  ND2CHD U80 ( .I1(n109), .I2(n110), .O(n447) );
  AOI222BHD U81 ( .A1(P[40]), .A2(n81), .B1(N132), .B2(n74), .C1(n62), .C2(
        X5x[0]), .O(n110) );
  AOI22BHD U82 ( .A1(X4x[0]), .A2(n88), .B1(N429), .B2(n69), .O(n109) );
  OAI112BHD U83 ( .C1(n113), .C2(n114), .A1(n115), .B1(n116), .O(n446) );
  AOI222BHD U84 ( .A1(N83), .A2(n117), .B1(n88), .B2(n118), .C1(N75), .C2(n119), .O(n116) );
  ND2CHD U85 ( .I1(n72), .I2(X5x[0]), .O(n115) );
  INVCHD U86 ( .I(X4x[0]), .O(n114) );
  OAI112BHD U87 ( .C1(n113), .C2(n120), .A1(n121), .B1(n122), .O(n445) );
  AOI222BHD U88 ( .A1(N84), .A2(n117), .B1(n89), .B2(n123), .C1(N76), .C2(n119), .O(n122) );
  ND2CHD U89 ( .I1(n72), .I2(X5x[1]), .O(n121) );
  INVCHD U90 ( .I(X4x[1]), .O(n120) );
  OAI112BHD U91 ( .C1(n113), .C2(n124), .A1(n125), .B1(n126), .O(n444) );
  AOI222BHD U92 ( .A1(N85), .A2(n117), .B1(n90), .B2(n127), .C1(N77), .C2(n119), .O(n126) );
  ND2CHD U93 ( .I1(n72), .I2(X5x[2]), .O(n125) );
  INVCHD U94 ( .I(X4x[2]), .O(n124) );
  OAI112BHD U95 ( .C1(n113), .C2(n128), .A1(n129), .B1(n130), .O(n443) );
  AOI222BHD U96 ( .A1(N86), .A2(n117), .B1(n90), .B2(n131), .C1(N78), .C2(n119), .O(n130) );
  ND2CHD U97 ( .I1(n71), .I2(X5x[3]), .O(n129) );
  INVCHD U98 ( .I(X4x[3]), .O(n128) );
  OAI112BHD U99 ( .C1(n113), .C2(n132), .A1(n133), .B1(n134), .O(n442) );
  AOI222BHD U100 ( .A1(N87), .A2(n117), .B1(n89), .B2(n135), .C1(N79), .C2(
        n119), .O(n134) );
  ND2CHD U101 ( .I1(n72), .I2(X5x[4]), .O(n133) );
  INVCHD U102 ( .I(X4x[4]), .O(n132) );
  OAI112BHD U103 ( .C1(n113), .C2(n136), .A1(n137), .B1(n138), .O(n441) );
  AOI222BHD U104 ( .A1(N88), .A2(n117), .B1(n89), .B2(n139), .C1(N80), .C2(
        n119), .O(n138) );
  ND2CHD U105 ( .I1(n72), .I2(X5x[5]), .O(n137) );
  INVCHD U106 ( .I(X4x[5]), .O(n136) );
  OAI112BHD U107 ( .C1(n113), .C2(n140), .A1(n141), .B1(n142), .O(n440) );
  AOI222BHD U108 ( .A1(N89), .A2(n117), .B1(n89), .B2(n143), .C1(N81), .C2(
        n119), .O(n142) );
  ND2CHD U109 ( .I1(n71), .I2(X5x[6]), .O(n141) );
  INVCHD U110 ( .I(X4x[6]), .O(n140) );
  OAI112BHD U111 ( .C1(n113), .C2(n144), .A1(n145), .B1(n146), .O(n439) );
  AOI222BHD U112 ( .A1(N90), .A2(n117), .B1(n90), .B2(n147), .C1(N82), .C2(
        n119), .O(n146) );
  ND2CHD U113 ( .I1(n72), .I2(X5x[7]), .O(n145) );
  INVCHD U114 ( .I(X4x[7]), .O(n144) );
  ND2CHD U115 ( .I1(n148), .I2(n149), .O(n438) );
  AOI222BHD U116 ( .A1(P[41]), .A2(n80), .B1(N133), .B2(n74), .C1(n62), .C2(
        X5x[1]), .O(n149) );
  AOI22BHD U117 ( .A1(X4x[1]), .A2(n88), .B1(N430), .B2(n69), .O(n148) );
  ND2CHD U118 ( .I1(n150), .I2(n151), .O(n437) );
  AOI222BHD U119 ( .A1(P[42]), .A2(n80), .B1(N134), .B2(n74), .C1(n62), .C2(
        X5x[2]), .O(n151) );
  AOI22BHD U120 ( .A1(X4x[2]), .A2(n88), .B1(N431), .B2(n68), .O(n150) );
  ND2CHD U121 ( .I1(n152), .I2(n153), .O(n436) );
  AOI222BHD U122 ( .A1(P[43]), .A2(n80), .B1(N135), .B2(n74), .C1(n62), .C2(
        X5x[3]), .O(n153) );
  AOI22BHD U123 ( .A1(X4x[3]), .A2(n88), .B1(N432), .B2(n70), .O(n152) );
  ND2CHD U124 ( .I1(n154), .I2(n155), .O(n435) );
  AOI222BHD U125 ( .A1(P[44]), .A2(n80), .B1(N136), .B2(n74), .C1(n62), .C2(
        X5x[4]), .O(n155) );
  AOI22BHD U126 ( .A1(X4x[4]), .A2(n88), .B1(N433), .B2(n70), .O(n154) );
  ND2CHD U127 ( .I1(n156), .I2(n157), .O(n434) );
  AOI222BHD U128 ( .A1(P[45]), .A2(n80), .B1(N137), .B2(n74), .C1(n62), .C2(
        X5x[5]), .O(n157) );
  AOI22BHD U129 ( .A1(X4x[5]), .A2(n88), .B1(N434), .B2(n69), .O(n156) );
  ND2CHD U130 ( .I1(n158), .I2(n159), .O(n433) );
  AOI222BHD U131 ( .A1(P[46]), .A2(n80), .B1(N138), .B2(n74), .C1(n62), .C2(
        X5x[6]), .O(n159) );
  AOI22BHD U132 ( .A1(X4x[6]), .A2(n88), .B1(N435), .B2(n69), .O(n158) );
  ND2CHD U133 ( .I1(n160), .I2(n161), .O(n432) );
  AOI222BHD U134 ( .A1(P[47]), .A2(n80), .B1(N139), .B2(n74), .C1(n62), .C2(
        X5x[7]), .O(n161) );
  AOI22BHD U135 ( .A1(X4x[7]), .A2(n89), .B1(N436), .B2(n70), .O(n160) );
  AO2222BHD U136 ( .A1(X7x[0]), .A2(n72), .B1(N197), .B2(n93), .C1(n63), .C2(
        X6x[0]), .D1(n84), .D2(n163), .O(n431) );
  XOR2CHD U137 ( .I1(WK3_7[0]), .I2(P[48]), .O(n163) );
  AO2222BHD U138 ( .A1(X7x[1]), .A2(n73), .B1(N198), .B2(n92), .C1(n63), .C2(
        X6x[1]), .D1(n83), .D2(n164), .O(n430) );
  XOR2CHD U139 ( .I1(WK3_7[1]), .I2(P[49]), .O(n164) );
  AO2222BHD U140 ( .A1(X7x[2]), .A2(n72), .B1(N199), .B2(n93), .C1(n63), .C2(
        X6x[2]), .D1(n84), .D2(n165), .O(n429) );
  XOR2CHD U141 ( .I1(WK3_7[2]), .I2(P[50]), .O(n165) );
  AO2222BHD U142 ( .A1(X7x[3]), .A2(n72), .B1(N200), .B2(n92), .C1(n63), .C2(
        X6x[3]), .D1(n83), .D2(n166), .O(n428) );
  XOR2CHD U143 ( .I1(WK3_7[3]), .I2(P[51]), .O(n166) );
  AO2222BHD U144 ( .A1(X7x[4]), .A2(n72), .B1(N201), .B2(n92), .C1(n63), .C2(
        X6x[4]), .D1(n84), .D2(n167), .O(n427) );
  XOR2CHD U145 ( .I1(WK3_7[4]), .I2(P[52]), .O(n167) );
  AO2222BHD U146 ( .A1(X7x[5]), .A2(n73), .B1(N202), .B2(n93), .C1(n63), .C2(
        X6x[5]), .D1(n83), .D2(n168), .O(n426) );
  XOR2CHD U147 ( .I1(WK3_7[5]), .I2(P[53]), .O(n168) );
  AO2222BHD U148 ( .A1(X7x[6]), .A2(n72), .B1(N203), .B2(n92), .C1(n63), .C2(
        X6x[6]), .D1(n83), .D2(n169), .O(n425) );
  XOR2CHD U149 ( .I1(WK3_7[6]), .I2(P[54]), .O(n169) );
  AO2222BHD U150 ( .A1(X7x[7]), .A2(n73), .B1(N204), .B2(n92), .C1(n63), .C2(
        X6x[7]), .D1(n84), .D2(n170), .O(n424) );
  XOR2CHD U151 ( .I1(WK3_7[7]), .I2(P[55]), .O(n170) );
  OAI112BHD U152 ( .C1(n179), .C2(n180), .A1(n181), .B1(n183), .O(n423) );
  AOI22BHD U153 ( .A1(P[56]), .A2(n82), .B1(n91), .B2(X6x[0]), .O(n183) );
  AOI22BHD U154 ( .A1(n184), .A2(n68), .B1(n185), .B2(n76), .O(n181) );
  XOR2CHD U155 ( .I1(X00x[0]), .I2(N437), .O(n184) );
  INVCHD U156 ( .I(X7x[0]), .O(n180) );
  OAI112BHD U157 ( .C1(n179), .C2(n186), .A1(n187), .B1(n188), .O(n422) );
  AOI22BHD U158 ( .A1(P[57]), .A2(n82), .B1(n91), .B2(X6x[1]), .O(n188) );
  AOI22BHD U159 ( .A1(n189), .A2(n68), .B1(n190), .B2(n76), .O(n187) );
  XOR2CHD U160 ( .I1(X00x[1]), .I2(N438), .O(n189) );
  INVCHD U161 ( .I(X7x[1]), .O(n186) );
  OAI112BHD U162 ( .C1(n179), .C2(n191), .A1(n192), .B1(n193), .O(n421) );
  AOI22BHD U163 ( .A1(P[58]), .A2(n81), .B1(n91), .B2(X6x[2]), .O(n193) );
  AOI22BHD U164 ( .A1(n194), .A2(n68), .B1(n195), .B2(n76), .O(n192) );
  XOR2CHD U165 ( .I1(X00x[2]), .I2(N439), .O(n194) );
  INVCHD U166 ( .I(X7x[2]), .O(n191) );
  OAI112BHD U167 ( .C1(n179), .C2(n196), .A1(n197), .B1(n198), .O(n420) );
  AOI22BHD U168 ( .A1(P[59]), .A2(n82), .B1(n91), .B2(X6x[3]), .O(n198) );
  AOI22BHD U169 ( .A1(n199), .A2(n68), .B1(n200), .B2(n76), .O(n197) );
  XOR2CHD U170 ( .I1(X00x[3]), .I2(N440), .O(n199) );
  INVCHD U171 ( .I(X7x[3]), .O(n196) );
  OAI112BHD U172 ( .C1(n179), .C2(n201), .A1(n202), .B1(n203), .O(n419) );
  AOI22BHD U173 ( .A1(P[60]), .A2(n81), .B1(n91), .B2(X6x[4]), .O(n203) );
  AOI22BHD U174 ( .A1(n204), .A2(n68), .B1(n205), .B2(n76), .O(n202) );
  XOR2CHD U175 ( .I1(X00x[4]), .I2(N441), .O(n204) );
  INVCHD U176 ( .I(X7x[4]), .O(n201) );
  OAI112BHD U177 ( .C1(n179), .C2(n206), .A1(n207), .B1(n208), .O(n418) );
  AOI22BHD U178 ( .A1(P[61]), .A2(n82), .B1(n91), .B2(X6x[5]), .O(n208) );
  AOI22BHD U179 ( .A1(n209), .A2(n68), .B1(n210), .B2(n76), .O(n207) );
  XOR2CHD U180 ( .I1(X00x[5]), .I2(N442), .O(n209) );
  INVCHD U181 ( .I(X7x[5]), .O(n206) );
  OAI112BHD U182 ( .C1(n179), .C2(n211), .A1(n212), .B1(n213), .O(n417) );
  AOI22BHD U183 ( .A1(P[62]), .A2(n81), .B1(n91), .B2(X6x[6]), .O(n213) );
  AOI22BHD U184 ( .A1(n214), .A2(n68), .B1(n215), .B2(n76), .O(n212) );
  XOR2CHD U185 ( .I1(X00x[6]), .I2(N443), .O(n214) );
  INVCHD U186 ( .I(X7x[6]), .O(n211) );
  OAI112BHD U187 ( .C1(n179), .C2(n216), .A1(n217), .B1(n218), .O(n416) );
  AOI22BHD U188 ( .A1(P[63]), .A2(n81), .B1(n91), .B2(X6x[7]), .O(n218) );
  AOI22BHD U189 ( .A1(n219), .A2(n68), .B1(n220), .B2(n76), .O(n217) );
  XOR2CHD U190 ( .I1(X00x[7]), .I2(N444), .O(n219) );
  INVCHD U191 ( .I(X7x[7]), .O(n216) );
  OAI112BHD U192 ( .C1(n113), .C2(n221), .A1(n222), .B1(n223), .O(n415) );
  AOI222BHD U193 ( .A1(N51), .A2(n117), .B1(n90), .B2(n185), .C1(N43), .C2(
        n119), .O(n223) );
  XOR2CHD U194 ( .I1(X7x[0]), .I2(N140), .O(n185) );
  ND2CHD U195 ( .I1(X1x[0]), .I2(n69), .O(n222) );
  INVCHD U196 ( .I(X0x[0]), .O(n221) );
  OAI112BHD U197 ( .C1(n113), .C2(n224), .A1(n225), .B1(n226), .O(n414) );
  AOI222BHD U198 ( .A1(N52), .A2(n117), .B1(n89), .B2(n190), .C1(N44), .C2(
        n119), .O(n226) );
  XOR2CHD U199 ( .I1(X7x[1]), .I2(N141), .O(n190) );
  ND2CHD U200 ( .I1(X1x[1]), .I2(n69), .O(n225) );
  INVCHD U201 ( .I(X0x[1]), .O(n224) );
  OAI112BHD U202 ( .C1(n113), .C2(n227), .A1(n228), .B1(n229), .O(n413) );
  AOI222BHD U203 ( .A1(N53), .A2(n117), .B1(n90), .B2(n195), .C1(N45), .C2(
        n119), .O(n229) );
  XOR2CHD U204 ( .I1(X7x[2]), .I2(N142), .O(n195) );
  ND2CHD U205 ( .I1(X1x[2]), .I2(n69), .O(n228) );
  INVCHD U206 ( .I(X0x[2]), .O(n227) );
  OAI112BHD U207 ( .C1(n113), .C2(n230), .A1(n231), .B1(n232), .O(n412) );
  AOI222BHD U208 ( .A1(N54), .A2(n117), .B1(n90), .B2(n200), .C1(N46), .C2(
        n119), .O(n232) );
  XOR2CHD U209 ( .I1(X7x[3]), .I2(N143), .O(n200) );
  ND2CHD U210 ( .I1(X1x[3]), .I2(n69), .O(n231) );
  INVCHD U211 ( .I(X0x[3]), .O(n230) );
  OAI112BHD U212 ( .C1(n113), .C2(n233), .A1(n234), .B1(n235), .O(n411) );
  AOI222BHD U213 ( .A1(N55), .A2(n117), .B1(n90), .B2(n205), .C1(N47), .C2(
        n119), .O(n235) );
  XOR2CHD U214 ( .I1(X7x[4]), .I2(N144), .O(n205) );
  ND2CHD U215 ( .I1(X1x[4]), .I2(n69), .O(n234) );
  INVCHD U216 ( .I(X0x[4]), .O(n233) );
  OAI112BHD U217 ( .C1(n113), .C2(n236), .A1(n237), .B1(n238), .O(n410) );
  AOI222BHD U218 ( .A1(N56), .A2(n117), .B1(n90), .B2(n210), .C1(N48), .C2(
        n119), .O(n238) );
  XOR2CHD U219 ( .I1(X7x[5]), .I2(N145), .O(n210) );
  ND2CHD U220 ( .I1(X1x[5]), .I2(n68), .O(n237) );
  INVCHD U221 ( .I(X0x[5]), .O(n236) );
  OAI112BHD U222 ( .C1(n113), .C2(n239), .A1(n240), .B1(n241), .O(n409) );
  AOI222BHD U223 ( .A1(N57), .A2(n117), .B1(n90), .B2(n215), .C1(N49), .C2(
        n119), .O(n241) );
  XOR2CHD U224 ( .I1(X7x[6]), .I2(N146), .O(n215) );
  ND2CHD U225 ( .I1(X1x[6]), .I2(n69), .O(n240) );
  INVCHD U226 ( .I(X0x[6]), .O(n239) );
  OAI112BHD U227 ( .C1(n113), .C2(n242), .A1(n243), .B1(n244), .O(n408) );
  AOI222BHD U228 ( .A1(N58), .A2(n117), .B1(n90), .B2(n220), .C1(N50), .C2(
        n119), .O(n244) );
  XOR2CHD U229 ( .I1(X7x[7]), .I2(N147), .O(n220) );
  ND2CHD U230 ( .I1(X1x[7]), .I2(n68), .O(n243) );
  INVCHD U231 ( .I(X0x[7]), .O(n242) );
  AO222CHD U232 ( .A1(N255), .A2(n247), .B1(N263), .B2(n64), .C1(C[0]), .C2(
        n103), .O(n407) );
  AO222CHD U233 ( .A1(N256), .A2(n247), .B1(N264), .B2(n64), .C1(C[1]), .C2(
        n103), .O(n406) );
  AO222CHD U234 ( .A1(N257), .A2(n247), .B1(N265), .B2(n64), .C1(C[2]), .C2(
        n103), .O(n405) );
  AO222CHD U235 ( .A1(N258), .A2(n247), .B1(N266), .B2(n64), .C1(C[3]), .C2(
        n103), .O(n404) );
  AO222CHD U236 ( .A1(N259), .A2(n247), .B1(N267), .B2(n64), .C1(C[4]), .C2(
        n103), .O(n403) );
  AO222CHD U237 ( .A1(N260), .A2(n247), .B1(N268), .B2(n64), .C1(C[5]), .C2(
        n103), .O(n402) );
  AO222CHD U238 ( .A1(N261), .A2(n247), .B1(N269), .B2(n64), .C1(C[6]), .C2(
        n103), .O(n401) );
  AO222CHD U239 ( .A1(N262), .A2(n247), .B1(N270), .B2(n64), .C1(C[7]), .C2(
        n103), .O(n400) );
  ND2CHD U240 ( .I1(n249), .I2(n250), .O(n399) );
  AOI222BHD U241 ( .A1(P[8]), .A2(n80), .B1(N108), .B2(n75), .C1(X1x[0]), .C2(
        n62), .O(n250) );
  AOI22BHD U242 ( .A1(X0x[0]), .A2(n89), .B1(N397), .B2(n70), .O(n249) );
  ND2CHD U243 ( .I1(n251), .I2(n252), .O(n398) );
  AOI222BHD U244 ( .A1(P[9]), .A2(n80), .B1(N109), .B2(n74), .C1(X1x[1]), .C2(
        n62), .O(n252) );
  AOI22BHD U245 ( .A1(X0x[1]), .A2(n89), .B1(N398), .B2(n70), .O(n251) );
  ND2CHD U246 ( .I1(n253), .I2(n254), .O(n397) );
  AOI222BHD U247 ( .A1(P[10]), .A2(n80), .B1(N110), .B2(n75), .C1(X1x[2]), 
        .C2(n62), .O(n254) );
  AOI22BHD U248 ( .A1(X0x[2]), .A2(n88), .B1(N399), .B2(n70), .O(n253) );
  ND2CHD U249 ( .I1(n255), .I2(n256), .O(n396) );
  AOI222BHD U250 ( .A1(P[11]), .A2(n80), .B1(N111), .B2(n75), .C1(X1x[3]), 
        .C2(n62), .O(n256) );
  AOI22BHD U251 ( .A1(X0x[3]), .A2(n89), .B1(N400), .B2(n70), .O(n255) );
  ND2CHD U252 ( .I1(n257), .I2(n258), .O(n395) );
  AOI222BHD U253 ( .A1(P[12]), .A2(n81), .B1(N112), .B2(n75), .C1(X1x[4]), 
        .C2(n62), .O(n258) );
  AOI22BHD U254 ( .A1(X0x[4]), .A2(n89), .B1(N401), .B2(n70), .O(n257) );
  ND2CHD U255 ( .I1(n259), .I2(n260), .O(n394) );
  AOI222BHD U256 ( .A1(P[13]), .A2(n81), .B1(N113), .B2(n74), .C1(X1x[5]), 
        .C2(n62), .O(n260) );
  AOI22BHD U257 ( .A1(X0x[5]), .A2(n88), .B1(N402), .B2(n70), .O(n259) );
  ND2CHD U258 ( .I1(n261), .I2(n262), .O(n393) );
  AOI222BHD U259 ( .A1(P[14]), .A2(n81), .B1(N114), .B2(n75), .C1(X1x[6]), 
        .C2(n62), .O(n262) );
  AOI22BHD U260 ( .A1(X0x[6]), .A2(n89), .B1(N403), .B2(n70), .O(n261) );
  ND2CHD U261 ( .I1(n263), .I2(n264), .O(n392) );
  AOI222BHD U262 ( .A1(P[15]), .A2(n81), .B1(N115), .B2(n74), .C1(X1x[7]), 
        .C2(n62), .O(n264) );
  AOI22BHD U263 ( .A1(X0x[7]), .A2(n88), .B1(N404), .B2(n69), .O(n263) );
  AO2222BHD U264 ( .A1(X3x[0]), .A2(n73), .B1(N173), .B2(n92), .C1(n63), .C2(
        X2x[0]), .D1(n83), .D2(n265), .O(n391) );
  XOR2CHD U265 ( .I1(WK1_5[0]), .I2(P[16]), .O(n265) );
  AO2222BHD U266 ( .A1(X3x[1]), .A2(n73), .B1(N174), .B2(n93), .C1(n63), .C2(
        X2x[1]), .D1(n83), .D2(n266), .O(n390) );
  XOR2CHD U267 ( .I1(WK1_5[1]), .I2(P[17]), .O(n266) );
  AO2222BHD U268 ( .A1(X3x[2]), .A2(n73), .B1(N175), .B2(n93), .C1(n63), .C2(
        X2x[2]), .D1(n83), .D2(n267), .O(n389) );
  XOR2CHD U269 ( .I1(WK1_5[2]), .I2(P[18]), .O(n267) );
  AO2222BHD U270 ( .A1(X3x[3]), .A2(n73), .B1(N176), .B2(n93), .C1(n63), .C2(
        X2x[3]), .D1(n83), .D2(n268), .O(n388) );
  XOR2CHD U271 ( .I1(WK1_5[3]), .I2(P[19]), .O(n268) );
  AO2222BHD U272 ( .A1(X3x[4]), .A2(n73), .B1(N177), .B2(n93), .C1(n63), .C2(
        X2x[4]), .D1(n83), .D2(n269), .O(n387) );
  XOR2CHD U273 ( .I1(WK1_5[4]), .I2(P[20]), .O(n269) );
  AO2222BHD U274 ( .A1(X3x[5]), .A2(n73), .B1(N178), .B2(n93), .C1(n63), .C2(
        X2x[5]), .D1(n83), .D2(n270), .O(n386) );
  XOR2CHD U275 ( .I1(WK1_5[5]), .I2(P[21]), .O(n270) );
  AO2222BHD U276 ( .A1(X3x[6]), .A2(n73), .B1(N179), .B2(n93), .C1(n63), .C2(
        X2x[6]), .D1(n83), .D2(n271), .O(n385) );
  XOR2CHD U277 ( .I1(WK1_5[6]), .I2(P[22]), .O(n271) );
  AO2222BHD U278 ( .A1(X3x[7]), .A2(n73), .B1(N180), .B2(n93), .C1(n63), .C2(
        X2x[7]), .D1(n83), .D2(n272), .O(n384) );
  XOR2CHD U279 ( .I1(WK1_5[7]), .I2(P[23]), .O(n272) );
  OAI112BHD U280 ( .C1(n179), .C2(n273), .A1(n274), .B1(n275), .O(n383) );
  AOI22BHD U281 ( .A1(P[24]), .A2(n81), .B1(n92), .B2(X2x[0]), .O(n275) );
  AOI22BHD U282 ( .A1(n71), .A2(n276), .B1(n118), .B2(n76), .O(n274) );
  XOR2CHD U283 ( .I1(X3x[0]), .I2(N116), .O(n118) );
  XOR2CHD U284 ( .I1(X4x[0]), .I2(N405), .O(n276) );
  INVCHD U285 ( .I(X3x[0]), .O(n273) );
  OAI112BHD U286 ( .C1(n179), .C2(n277), .A1(n278), .B1(n279), .O(n382) );
  AOI22BHD U287 ( .A1(P[25]), .A2(n82), .B1(n91), .B2(X2x[1]), .O(n279) );
  AOI22BHD U288 ( .A1(n71), .A2(n280), .B1(n123), .B2(n75), .O(n278) );
  XOR2CHD U289 ( .I1(X3x[1]), .I2(N117), .O(n123) );
  XOR2CHD U290 ( .I1(X4x[1]), .I2(N406), .O(n280) );
  INVCHD U291 ( .I(X3x[1]), .O(n277) );
  OAI112BHD U292 ( .C1(n179), .C2(n281), .A1(n282), .B1(n283), .O(n381) );
  AOI22BHD U293 ( .A1(P[26]), .A2(n81), .B1(n91), .B2(X2x[2]), .O(n283) );
  AOI22BHD U294 ( .A1(n71), .A2(n284), .B1(n127), .B2(n75), .O(n282) );
  XOR2CHD U295 ( .I1(X3x[2]), .I2(N118), .O(n127) );
  XOR2CHD U296 ( .I1(X4x[2]), .I2(N407), .O(n284) );
  INVCHD U297 ( .I(X3x[2]), .O(n281) );
  OAI112BHD U298 ( .C1(n179), .C2(n285), .A1(n286), .B1(n287), .O(n380) );
  AOI22BHD U299 ( .A1(P[27]), .A2(n82), .B1(n92), .B2(X2x[3]), .O(n287) );
  AOI22BHD U300 ( .A1(n71), .A2(n288), .B1(n131), .B2(n76), .O(n286) );
  XOR2CHD U301 ( .I1(X3x[3]), .I2(N119), .O(n131) );
  XOR2CHD U302 ( .I1(X4x[3]), .I2(N408), .O(n288) );
  INVCHD U303 ( .I(X3x[3]), .O(n285) );
  OAI112BHD U304 ( .C1(n179), .C2(n289), .A1(n290), .B1(n291), .O(n379) );
  AOI22BHD U305 ( .A1(P[28]), .A2(n82), .B1(n92), .B2(X2x[4]), .O(n291) );
  AOI22BHD U306 ( .A1(n71), .A2(n292), .B1(n135), .B2(n75), .O(n290) );
  XOR2CHD U307 ( .I1(X3x[4]), .I2(N120), .O(n135) );
  XOR2CHD U308 ( .I1(X4x[4]), .I2(N409), .O(n292) );
  INVCHD U309 ( .I(X3x[4]), .O(n289) );
  OAI112BHD U310 ( .C1(n179), .C2(n293), .A1(n294), .B1(n295), .O(n378) );
  AOI22BHD U311 ( .A1(P[29]), .A2(n82), .B1(n91), .B2(X2x[5]), .O(n295) );
  AOI22BHD U312 ( .A1(n71), .A2(n296), .B1(n139), .B2(n75), .O(n294) );
  XOR2CHD U313 ( .I1(X3x[5]), .I2(N121), .O(n139) );
  XOR2CHD U314 ( .I1(X4x[5]), .I2(N410), .O(n296) );
  INVCHD U315 ( .I(X3x[5]), .O(n293) );
  OAI112BHD U316 ( .C1(n179), .C2(n297), .A1(n298), .B1(n299), .O(n377) );
  AOI22BHD U317 ( .A1(P[30]), .A2(n82), .B1(n92), .B2(X2x[6]), .O(n299) );
  AOI22BHD U318 ( .A1(n71), .A2(n300), .B1(n143), .B2(n75), .O(n298) );
  XOR2CHD U319 ( .I1(X3x[6]), .I2(N122), .O(n143) );
  XOR2CHD U320 ( .I1(X4x[6]), .I2(N411), .O(n300) );
  INVCHD U321 ( .I(X3x[6]), .O(n297) );
  OAI112BHD U322 ( .C1(n179), .C2(n301), .A1(n302), .B1(n303), .O(n376) );
  AOI22BHD U323 ( .A1(P[31]), .A2(n82), .B1(n92), .B2(X2x[7]), .O(n303) );
  AOI22BHD U324 ( .A1(n70), .A2(n304), .B1(n147), .B2(n75), .O(n302) );
  XOR2CHD U325 ( .I1(X3x[7]), .I2(N123), .O(n147) );
  XOR2CHD U326 ( .I1(X4x[7]), .I2(N412), .O(n304) );
  INVCHD U327 ( .I(X3x[7]), .O(n301) );
  INVCHD U328 ( .I(n245), .O(n111) );
  ND3CHD U329 ( .I1(n108), .I2(n306), .I3(n307), .O(n245) );
  OR2B1CHD U330 ( .I1(n310), .B1(n108), .O(n308) );
  XOR2CHD U331 ( .I1(n108), .I2(n307), .O(n309) );
  NR2BHD U332 ( .I1(n311), .I2(n310), .O(n307) );
  AO222CHD U333 ( .A1(N294), .A2(n247), .B1(N302), .B2(n64), .C1(C[39]), .C2(
        n102), .O(n375) );
  AO222CHD U334 ( .A1(N293), .A2(n247), .B1(N301), .B2(n64), .C1(C[38]), .C2(
        n102), .O(n374) );
  AO222CHD U335 ( .A1(N292), .A2(n247), .B1(N300), .B2(n64), .C1(C[37]), .C2(
        n102), .O(n373) );
  AO222CHD U336 ( .A1(N291), .A2(n247), .B1(N299), .B2(n64), .C1(C[36]), .C2(
        n102), .O(n372) );
  AO222CHD U337 ( .A1(N290), .A2(n247), .B1(N298), .B2(n64), .C1(C[35]), .C2(
        n102), .O(n371) );
  AO222CHD U338 ( .A1(N289), .A2(n247), .B1(N297), .B2(n64), .C1(C[34]), .C2(
        n102), .O(n370) );
  AO222CHD U339 ( .A1(N288), .A2(n247), .B1(N296), .B2(n64), .C1(C[33]), .C2(
        n102), .O(n369) );
  AO222CHD U340 ( .A1(N287), .A2(n247), .B1(N295), .B2(n64), .C1(C[32]), .C2(
        n102), .O(n368) );
  INVCHD U341 ( .I(ed), .O(n246) );
  ND2CHD U342 ( .I1(n305), .I2(i_round[5]), .O(n182) );
  NR3BHD U343 ( .I1(n310), .I2(n107), .I3(n306), .O(n305) );
  XOR4EHD U344 ( .I1(X0x[0]), .I2(SKx0[4]), .I3(X0x[6]), .I4(X0x[1]), .O(N9)
         );
  XOR4EHD U345 ( .I1(X0x[1]), .I2(SKx0[5]), .I3(X0x[7]), .I4(X0x[2]), .O(N8)
         );
  XOR4EHD U346 ( .I1(X0x[0]), .I2(SKx0[6]), .I3(X0x[3]), .I4(X0x[2]), .O(N7)
         );
  XOR4EHD U347 ( .I1(X0x[1]), .I2(SKx0[7]), .I3(X0x[4]), .I4(X0x[3]), .O(N6)
         );
  XOR4EHD U348 ( .I1(n176), .I2(X5x[4]), .I3(SKx2[0]), .I4(n173), .O(N428) );
  XOR4EHD U349 ( .I1(n175), .I2(X5x[5]), .I3(SKx2[1]), .I4(n172), .O(N427) );
  XOR4EHD U350 ( .I1(n174), .I2(X5x[6]), .I3(SKx2[2]), .I4(n171), .O(N426) );
  XOR4EHD U351 ( .I1(n178), .I2(X5x[5]), .I3(SKx2[3]), .I4(n171), .O(N425) );
  XOR4EHD U352 ( .I1(n178), .I2(X5x[1]), .I3(SKx2[4]), .I4(n172), .O(N424) );
  XOR4EHD U353 ( .I1(n177), .I2(X5x[2]), .I3(SKx2[5]), .I4(n171), .O(N423) );
  XOR4EHD U354 ( .I1(n178), .I2(X5x[2]), .I3(SKx2[6]), .I4(n175), .O(N422) );
  XOR4EHD U355 ( .I1(n177), .I2(X5x[3]), .I3(SKx2[7]), .I4(n174), .O(N421) );
  XOR4EHD U356 ( .I1(X1x[2]), .I2(SKx0[0]), .I3(X1x[5]), .I4(X1x[4]), .O(N396)
         );
  XOR4EHD U357 ( .I1(X1x[3]), .I2(SKx0[1]), .I3(X1x[6]), .I4(X1x[5]), .O(N395)
         );
  XOR4EHD U358 ( .I1(X1x[4]), .I2(SKx0[2]), .I3(X1x[7]), .I4(X1x[6]), .O(N394)
         );
  XOR4EHD U359 ( .I1(X1x[0]), .I2(SKx0[3]), .I3(X1x[7]), .I4(X1x[5]), .O(N393)
         );
  XOR4EHD U360 ( .I1(X1x[0]), .I2(SKx0[4]), .I3(X1x[6]), .I4(X1x[1]), .O(N392)
         );
  XOR4EHD U361 ( .I1(X1x[1]), .I2(SKx0[5]), .I3(X1x[7]), .I4(X1x[2]), .O(N391)
         );
  XOR4EHD U362 ( .I1(X1x[0]), .I2(SKx0[6]), .I3(X1x[3]), .I4(X1x[2]), .O(N390)
         );
  XOR4EHD U363 ( .I1(X1x[1]), .I2(SKx0[7]), .I3(X1x[4]), .I4(X1x[3]), .O(N389)
         );
  OAI112BHD U364 ( .C1(n311), .C2(n312), .A1(n310), .B1(i_round[5]), .O(N23)
         );
  ND3CHD U365 ( .I1(n105), .I2(n104), .I3(n106), .O(n310) );
  ND2CHD U366 ( .I1(n105), .I2(n104), .O(n312) );
  XOR4EHD U367 ( .I1(X4x[2]), .I2(SKx2[0]), .I3(X4x[5]), .I4(X4x[4]), .O(N21)
         );
  XOR4EHD U368 ( .I1(X4x[3]), .I2(SKx2[1]), .I3(X4x[6]), .I4(X4x[5]), .O(N20)
         );
  XOR4EHD U369 ( .I1(X4x[4]), .I2(SKx2[2]), .I3(X4x[7]), .I4(X4x[6]), .O(N19)
         );
  XOR4EHD U370 ( .I1(X4x[0]), .I2(SKx2[3]), .I3(X4x[7]), .I4(X4x[5]), .O(N18)
         );
  XOR4EHD U371 ( .I1(X4x[0]), .I2(SKx2[4]), .I3(X4x[6]), .I4(X4x[1]), .O(N17)
         );
  XOR4EHD U372 ( .I1(X4x[1]), .I2(SKx2[5]), .I3(X4x[7]), .I4(X4x[2]), .O(N16)
         );
  XOR4EHD U373 ( .I1(X4x[0]), .I2(SKx2[6]), .I3(X4x[3]), .I4(X4x[2]), .O(N15)
         );
  XOR4EHD U374 ( .I1(X4x[1]), .I2(SKx2[7]), .I3(X4x[4]), .I4(X4x[3]), .O(N14)
         );
  XOR4EHD U375 ( .I1(X0x[2]), .I2(SKx0[0]), .I3(X0x[5]), .I4(X0x[4]), .O(N13)
         );
  XOR4EHD U376 ( .I1(X0x[3]), .I2(SKx0[1]), .I3(X0x[6]), .I4(X0x[5]), .O(N12)
         );
  XOR4EHD U377 ( .I1(X0x[4]), .I2(SKx0[2]), .I3(X0x[7]), .I4(X0x[6]), .O(N11)
         );
  XOR4EHD U378 ( .I1(X0x[0]), .I2(SKx0[3]), .I3(X0x[7]), .I4(X0x[5]), .O(N10)
         );
  XOR3CHD U379 ( .I1(X7x[6]), .I2(X7x[5]), .I3(X7x[0]), .O(F0X7[7]) );
  XOR3CHD U380 ( .I1(X7x[7]), .I2(X7x[5]), .I3(X7x[4]), .O(F0X7[6]) );
  XOR3CHD U381 ( .I1(X7x[6]), .I2(X7x[4]), .I3(X7x[3]), .O(F0X7[5]) );
  XOR3CHD U382 ( .I1(X7x[5]), .I2(X7x[3]), .I3(X7x[2]), .O(F0X7[4]) );
  XOR3CHD U383 ( .I1(X7x[4]), .I2(X7x[2]), .I3(X7x[1]), .O(F0X7[3]) );
  XOR3CHD U384 ( .I1(X7x[3]), .I2(X7x[1]), .I3(X7x[0]), .O(F0X7[2]) );
  XOR3CHD U385 ( .I1(X7x[7]), .I2(X7x[2]), .I3(X7x[0]), .O(F0X7[1]) );
  XOR3CHD U386 ( .I1(X7x[7]), .I2(X7x[6]), .I3(X7x[1]), .O(F0X7[0]) );
  XOR3CHD U387 ( .I1(X6x[6]), .I2(X6x[5]), .I3(X6x[0]), .O(F0X6[7]) );
  XOR3CHD U388 ( .I1(X6x[7]), .I2(X6x[5]), .I3(X6x[4]), .O(F0X6[6]) );
  XOR3CHD U389 ( .I1(X6x[6]), .I2(X6x[4]), .I3(X6x[3]), .O(F0X6[5]) );
  XOR3CHD U390 ( .I1(X6x[5]), .I2(X6x[3]), .I3(X6x[2]), .O(F0X6[4]) );
  XOR3CHD U391 ( .I1(X6x[4]), .I2(X6x[2]), .I3(X6x[1]), .O(F0X6[3]) );
  XOR3CHD U392 ( .I1(X6x[3]), .I2(X6x[1]), .I3(X6x[0]), .O(F0X6[2]) );
  XOR3CHD U393 ( .I1(X6x[7]), .I2(X6x[2]), .I3(X6x[0]), .O(F0X6[1]) );
  XOR3CHD U394 ( .I1(X6x[7]), .I2(X6x[6]), .I3(X6x[1]), .O(F0X6[0]) );
  XOR3CHD U395 ( .I1(X3x[6]), .I2(X3x[5]), .I3(X3x[0]), .O(F0X3[7]) );
  XOR3CHD U396 ( .I1(X3x[5]), .I2(X3x[4]), .I3(X2x[7]), .O(F0X3[6]) );
  XOR3CHD U397 ( .I1(X3x[4]), .I2(X3x[3]), .I3(X2x[6]), .O(F0X3[5]) );
  XOR3CHD U398 ( .I1(X3x[3]), .I2(X3x[2]), .I3(X2x[5]), .O(F0X3[4]) );
  XOR3CHD U399 ( .I1(X3x[2]), .I2(X3x[1]), .I3(X2x[4]), .O(F0X3[3]) );
  XOR3CHD U400 ( .I1(X3x[1]), .I2(X3x[0]), .I3(X2x[3]), .O(F0X3[2]) );
  XOR2CHD U401 ( .I1(X3x[0]), .I2(n313), .O(F0X3[1]) );
  XOR2CHD U402 ( .I1(X3x[7]), .I2(n314), .O(F0X3[0]) );
  XOR3CHD U403 ( .I1(X2x[6]), .I2(X2x[5]), .I3(X2x[0]), .O(F0X2[7]) );
  XOR3CHD U404 ( .I1(X2x[7]), .I2(X2x[5]), .I3(X2x[4]), .O(F0X2[6]) );
  XOR3CHD U405 ( .I1(X2x[6]), .I2(X2x[4]), .I3(X2x[3]), .O(F0X2[5]) );
  XOR3CHD U406 ( .I1(X2x[5]), .I2(X2x[3]), .I3(X2x[2]), .O(F0X2[4]) );
  XOR3CHD U407 ( .I1(X2x[4]), .I2(X2x[2]), .I3(X2x[1]), .O(F0X2[3]) );
  XOR3CHD U408 ( .I1(X2x[3]), .I2(X2x[1]), .I3(X2x[0]), .O(F0X2[2]) );
  XOR2CHD U409 ( .I1(X2x[0]), .I2(n313), .O(F0X2[1]) );
  XOR2CHD U410 ( .I1(X2x[2]), .I2(X2x[7]), .O(n313) );
  XOR2CHD U411 ( .I1(X2x[7]), .I2(n314), .O(F0X2[0]) );
  XOR2CHD U412 ( .I1(X2x[1]), .I2(X2x[6]), .O(n314) );
endmodule


module SK_gen ( MK, clk, reset, ed, SKx0, SKx1, SKx2, SKx3 );
  input [127:0] MK;
  output [7:0] SKx0;
  output [7:0] SKx1;
  output [7:0] SKx2;
  output [7:0] SKx3;
  input clk, reset, ed;
  wire   N75, N76, N77, N78, N79, N89, N90, N91, N92, N93, n1, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543,
         \add_35/carry[5] , \add_35/carry[4] , \add_35/carry[3] ,
         \add_35/carry[2] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586;
  wire   [5:0] i_round;
  wire   [6:0] dx0;
  wire   [6:0] dx1;
  wire   [6:0] dx2;
  wire   [6:0] dx3;
  wire   [7:0] mkx0;
  wire   [7:0] mkx1;
  wire   [7:0] mkx2;
  wire   [7:0] mkx3;

  SK_gen_DW01_add_0 add_354 ( .A(mkx3), .B({n1, dx3}), .CI(n1), .SUM(SKx3) );
  SK_gen_DW01_add_1 add_353 ( .A(mkx2), .B({n1, dx2}), .CI(n1), .SUM(SKx2) );
  SK_gen_DW01_add_2 add_352 ( .A(mkx1), .B({n1, dx1}), .CI(n1), .SUM(SKx1) );
  SK_gen_DW01_add_3 add_351 ( .A(mkx0), .B({n1, dx0}), .CI(n1), .SUM(SKx0) );
  QDFFEHD \mkx0_reg[7]  ( .D(n509), .CK(clk), .Q(mkx0[7]) );
  QDFFEHD \mkx0_reg[6]  ( .D(n508), .CK(clk), .Q(mkx0[6]) );
  QDFFEHD \mkx0_reg[5]  ( .D(n507), .CK(clk), .Q(mkx0[5]) );
  QDFFEHD \mkx0_reg[4]  ( .D(n506), .CK(clk), .Q(mkx0[4]) );
  QDFFEHD \mkx0_reg[3]  ( .D(n505), .CK(clk), .Q(mkx0[3]) );
  QDFFEHD \mkx1_reg[7]  ( .D(n501), .CK(clk), .Q(mkx1[7]) );
  QDFFEHD \mkx1_reg[6]  ( .D(n500), .CK(clk), .Q(mkx1[6]) );
  QDFFEHD \mkx1_reg[5]  ( .D(n499), .CK(clk), .Q(mkx1[5]) );
  QDFFEHD \mkx1_reg[4]  ( .D(n498), .CK(clk), .Q(mkx1[4]) );
  QDFFEHD \mkx1_reg[3]  ( .D(n497), .CK(clk), .Q(mkx1[3]) );
  QDFFEHD \mkx1_reg[2]  ( .D(n496), .CK(clk), .Q(mkx1[2]) );
  QDFFEHD \mkx2_reg[7]  ( .D(n493), .CK(clk), .Q(mkx2[7]) );
  QDFFEHD \mkx2_reg[6]  ( .D(n492), .CK(clk), .Q(mkx2[6]) );
  QDFFEHD \mkx2_reg[5]  ( .D(n491), .CK(clk), .Q(mkx2[5]) );
  QDFFEHD \mkx2_reg[4]  ( .D(n490), .CK(clk), .Q(mkx2[4]) );
  QDFFEHD \mkx2_reg[3]  ( .D(n489), .CK(clk), .Q(mkx2[3]) );
  QDFFEHD \mkx3_reg[7]  ( .D(n485), .CK(clk), .Q(mkx3[7]) );
  QDFFEHD \mkx3_reg[6]  ( .D(n484), .CK(clk), .Q(mkx3[6]) );
  QDFFEHD \mkx3_reg[5]  ( .D(n483), .CK(clk), .Q(mkx3[5]) );
  QDFFEHD \mkx3_reg[4]  ( .D(n482), .CK(clk), .Q(mkx3[4]) );
  QDFFEHD \mkx3_reg[3]  ( .D(n481), .CK(clk), .Q(mkx3[3]) );
  QDFFEHD \mkx3_reg[2]  ( .D(n480), .CK(clk), .Q(mkx3[2]) );
  QDFFEHD \dx0_reg[6]  ( .D(n537), .CK(clk), .Q(dx0[6]) );
  QDFFEHD \dx0_reg[5]  ( .D(n536), .CK(clk), .Q(dx0[5]) );
  QDFFEHD \dx0_reg[4]  ( .D(n535), .CK(clk), .Q(dx0[4]) );
  QDFFEHD \dx0_reg[3]  ( .D(n534), .CK(clk), .Q(dx0[3]) );
  QDFFEHD \dx1_reg[6]  ( .D(n530), .CK(clk), .Q(dx1[6]) );
  QDFFEHD \dx1_reg[5]  ( .D(n529), .CK(clk), .Q(dx1[5]) );
  QDFFEHD \dx1_reg[4]  ( .D(n528), .CK(clk), .Q(dx1[4]) );
  QDFFEHD \dx1_reg[3]  ( .D(n527), .CK(clk), .Q(dx1[3]) );
  QDFFEHD \dx1_reg[2]  ( .D(n526), .CK(clk), .Q(dx1[2]) );
  QDFFEHD \dx2_reg[6]  ( .D(n523), .CK(clk), .Q(dx2[6]) );
  QDFFEHD \dx2_reg[5]  ( .D(n522), .CK(clk), .Q(dx2[5]) );
  QDFFEHD \dx2_reg[4]  ( .D(n521), .CK(clk), .Q(dx2[4]) );
  QDFFEHD \dx2_reg[3]  ( .D(n520), .CK(clk), .Q(dx2[3]) );
  QDFFEHD \dx3_reg[5]  ( .D(n515), .CK(clk), .Q(dx3[5]) );
  QDFFEHD \dx3_reg[4]  ( .D(n514), .CK(clk), .Q(dx3[4]) );
  QDFFEHD \dx3_reg[3]  ( .D(n513), .CK(clk), .Q(dx3[3]) );
  QDFFEHD \dx3_reg[2]  ( .D(n512), .CK(clk), .Q(dx3[2]) );
  QDFFEHD \dx3_reg[6]  ( .D(n516), .CK(clk), .Q(dx3[6]) );
  QDFFEHD \mkx0_reg[2]  ( .D(n504), .CK(clk), .Q(mkx0[2]) );
  QDFFEHD \mkx0_reg[1]  ( .D(n503), .CK(clk), .Q(mkx0[1]) );
  QDFFEHD \mkx0_reg[0]  ( .D(n502), .CK(clk), .Q(mkx0[0]) );
  QDFFEHD \mkx1_reg[1]  ( .D(n495), .CK(clk), .Q(mkx1[1]) );
  QDFFEHD \mkx1_reg[0]  ( .D(n494), .CK(clk), .Q(mkx1[0]) );
  QDFFEHD \mkx2_reg[2]  ( .D(n488), .CK(clk), .Q(mkx2[2]) );
  QDFFEHD \mkx2_reg[1]  ( .D(n487), .CK(clk), .Q(mkx2[1]) );
  QDFFEHD \mkx2_reg[0]  ( .D(n486), .CK(clk), .Q(mkx2[0]) );
  QDFFEHD \mkx3_reg[1]  ( .D(n479), .CK(clk), .Q(mkx3[1]) );
  QDFFEHD \mkx3_reg[0]  ( .D(n478), .CK(clk), .Q(mkx3[0]) );
  QDFFEHD \dx0_reg[2]  ( .D(n533), .CK(clk), .Q(dx0[2]) );
  QDFFEHD \dx0_reg[1]  ( .D(n532), .CK(clk), .Q(dx0[1]) );
  QDFFEHD \dx1_reg[1]  ( .D(n525), .CK(clk), .Q(dx1[1]) );
  QDFFEHD \dx1_reg[0]  ( .D(n524), .CK(clk), .Q(dx1[0]) );
  QDFFEHD \dx2_reg[2]  ( .D(n519), .CK(clk), .Q(dx2[2]) );
  QDFFEHD \dx2_reg[1]  ( .D(n518), .CK(clk), .Q(dx2[1]) );
  QDFFEHD \dx2_reg[0]  ( .D(n517), .CK(clk), .Q(dx2[0]) );
  QDFFEHD \dx3_reg[1]  ( .D(n511), .CK(clk), .Q(dx3[1]) );
  QDFFEHD \dx3_reg[0]  ( .D(n510), .CK(clk), .Q(dx3[0]) );
  QDFFEHD \dx0_reg[0]  ( .D(n531), .CK(clk), .Q(dx0[0]) );
  QDFFEHD \i_round_reg[3]  ( .D(n539), .CK(clk), .Q(i_round[3]) );
  QDFFEHD \i_round_reg[4]  ( .D(n538), .CK(clk), .Q(i_round[4]) );
  QDFFEHD \i_round_reg[5]  ( .D(n542), .CK(clk), .Q(i_round[5]) );
  QDFFEHD \i_round_reg[2]  ( .D(n540), .CK(clk), .Q(i_round[2]) );
  QDFFEHD \i_round_reg[0]  ( .D(n543), .CK(clk), .Q(i_round[0]) );
  QDFFEHD \i_round_reg[1]  ( .D(n541), .CK(clk), .Q(i_round[1]) );
  AOI12CHD U3 ( .B1(n124), .B2(n162), .A1(n115), .O(n2) );
  AOI12CHD U4 ( .B1(n582), .B2(n186), .A1(n153), .O(n3) );
  AOI12CHD U5 ( .B1(n131), .B2(n133), .A1(n152), .O(n4) );
  AOI12CHD U6 ( .B1(n162), .B2(n186), .A1(n140), .O(n5) );
  AOI12CHD U7 ( .B1(n133), .B2(n162), .A1(n158), .O(n6) );
  BUFEHD U8 ( .I(n71), .O(n69) );
  BUFEHD U9 ( .I(n72), .O(n68) );
  BUFEHD U10 ( .I(n72), .O(n67) );
  BUFEHD U11 ( .I(n71), .O(n70) );
  BUFEHD U12 ( .I(n206), .O(n71) );
  BUFEHD U13 ( .I(n206), .O(n72) );
  BUFEHD U14 ( .I(n21), .O(n24) );
  BUFEHD U15 ( .I(n21), .O(n23) );
  BUFEHD U16 ( .I(n22), .O(n25) );
  BUFEHD U17 ( .I(n22), .O(n26) );
  BUFEHD U18 ( .I(n30), .O(n32) );
  INVDHD U19 ( .I(n28), .O(n27) );
  INVDHD U20 ( .I(n11), .O(n9) );
  BUFEHD U21 ( .I(n8), .O(n11) );
  BUFEHD U22 ( .I(n54), .O(n53) );
  INVDHD U23 ( .I(n52), .O(n54) );
  BUFEHD U24 ( .I(n43), .O(n42) );
  INVDHD U25 ( .I(n113), .O(n121) );
  BUFEHD U26 ( .I(n14), .O(n13) );
  INVDHD U27 ( .I(n12), .O(n14) );
  INVDHD U28 ( .I(n58), .O(n55) );
  BUFEHD U29 ( .I(n60), .O(n58) );
  INVDHD U30 ( .I(n59), .O(n56) );
  BUFEHD U31 ( .I(n60), .O(n59) );
  BUFEHD U32 ( .I(n5), .O(n22) );
  BUFEHD U33 ( .I(n5), .O(n21) );
  BUFEHD U34 ( .I(n15), .O(n17) );
  BUFEHD U35 ( .I(n15), .O(n18) );
  BUFEHD U36 ( .I(n177), .O(n36) );
  BUFEHD U37 ( .I(n177), .O(n38) );
  BUFEHD U38 ( .I(n177), .O(n37) );
  BUFEHD U39 ( .I(n8), .O(n10) );
  BUFEHD U40 ( .I(n16), .O(n19) );
  BUFEHD U41 ( .I(n31), .O(n34) );
  BUFEHD U42 ( .I(n30), .O(n33) );
  BUFEHD U43 ( .I(n44), .O(n39) );
  BUFEHD U44 ( .I(n44), .O(n40) );
  BUFEHD U45 ( .I(n43), .O(n41) );
  BUFEHD U46 ( .I(n31), .O(n35) );
  BUFEHD U47 ( .I(n16), .O(n20) );
  BUFEHD U48 ( .I(n7), .O(n28) );
  BUFEHD U49 ( .I(n60), .O(n57) );
  INVDHD U50 ( .I(n189), .O(n60) );
  BUFEHD U51 ( .I(n188), .O(n52) );
  BUFEHD U52 ( .I(n45), .O(n43) );
  BUFEHD U53 ( .I(n4), .O(n30) );
  BUFEHD U54 ( .I(n3), .O(n51) );
  BUFEHD U55 ( .I(n2), .O(n48) );
  BUFEHD U56 ( .I(n143), .O(n12) );
  BUFEHD U57 ( .I(n7), .O(n29) );
  BUFEHD U58 ( .I(n6), .O(n16) );
  BUFEHD U59 ( .I(n6), .O(n15) );
  BUFEHD U60 ( .I(n45), .O(n44) );
  BUFEHD U61 ( .I(n4), .O(n31) );
  BUFEHD U62 ( .I(n2), .O(n46) );
  BUFEHD U63 ( .I(n2), .O(n47) );
  BUFEHD U64 ( .I(n3), .O(n49) );
  BUFEHD U65 ( .I(n3), .O(n50) );
  BUFEHD U66 ( .I(n65), .O(n63) );
  BUFEHD U67 ( .I(n66), .O(n62) );
  BUFEHD U68 ( .I(n66), .O(n61) );
  BUFEHD U69 ( .I(n65), .O(n64) );
  AOI12EHD U70 ( .B1(n142), .B2(n141), .A1(n159), .O(n118) );
  AN2EHD U71 ( .I1(n179), .I2(n180), .O(n94) );
  OA12EHD U72 ( .B1(n93), .B2(n145), .A1(n106), .O(n7) );
  AO12EHD U73 ( .B1(n142), .B2(n131), .A1(n170), .O(n8) );
  INVDHD U74 ( .I(n8), .O(n126) );
  BUFEHD U75 ( .I(n178), .O(n45) );
  INVDHD U76 ( .I(n73), .O(n77) );
  INVDHD U77 ( .I(n74), .O(n78) );
  BUFEHD U78 ( .I(n205), .O(n65) );
  BUFEHD U79 ( .I(n205), .O(n66) );
  NR2CHD U80 ( .I1(n583), .I2(i_round[1]), .O(n124) );
  HA1EHD U81 ( .A(i_round[1]), .B(i_round[0]), .C(\add_35/carry[2] ), .S(N75)
         );
  HA1EHD U82 ( .A(i_round[2]), .B(\add_35/carry[2] ), .C(\add_35/carry[3] ), 
        .S(N76) );
  HA1EHD U83 ( .A(i_round[3]), .B(\add_35/carry[3] ), .C(\add_35/carry[4] ), 
        .S(N77) );
  HA1EHD U84 ( .A(i_round[4]), .B(\add_35/carry[4] ), .C(\add_35/carry[5] ), 
        .S(N78) );
  TIE0DHD U85 ( .O(n1) );
  OA12EHD U86 ( .B1(n578), .B2(n145), .A1(n138), .O(n120) );
  XOR2CHD U87 ( .I1(\add_35/carry[5] ), .I2(i_round[5]), .O(N79) );
  NR2BHD U88 ( .I1(i_round[1]), .I2(i_round[0]), .O(n73) );
  AO12CHD U89 ( .B1(i_round[0]), .B2(i_round[1]), .A1(n73), .O(N89) );
  NR2BHD U90 ( .I1(n77), .I2(i_round[2]), .O(n74) );
  AO12CHD U91 ( .B1(n77), .B2(i_round[2]), .A1(n74), .O(N90) );
  NR2BHD U92 ( .I1(n78), .I2(i_round[3]), .O(n75) );
  AO12CHD U93 ( .B1(n78), .B2(i_round[3]), .A1(n75), .O(N91) );
  XOR2CHD U94 ( .I1(i_round[4]), .I2(n75), .O(N92) );
  AN2B1CHD U95 ( .I1(n75), .B1(i_round[4]), .O(n76) );
  XOR2CHD U96 ( .I1(i_round[5]), .I2(n76), .O(N93) );
  AO112CHD U97 ( .C1(n580), .C2(n79), .A1(n80), .B1(n81), .O(n543) );
  MUX2CHD U98 ( .A(n82), .B(n83), .S(i_round[0]), .O(n81) );
  OR3B2CHD U99 ( .I1(n80), .B1(n84), .B2(n85), .O(n542) );
  AOI22BHD U100 ( .A1(N93), .A2(n79), .B1(N79), .B2(n82), .O(n85) );
  NR2BHD U101 ( .I1(n86), .I2(ed), .O(n80) );
  AO222CHD U102 ( .A1(N89), .A2(n79), .B1(i_round[1]), .B2(n83), .C1(N75), 
        .C2(n82), .O(n541) );
  AO222CHD U103 ( .A1(N90), .A2(n79), .B1(i_round[2]), .B2(n83), .C1(N76), 
        .C2(n82), .O(n540) );
  AO222CHD U104 ( .A1(N91), .A2(n79), .B1(i_round[3]), .B2(n83), .C1(N77), 
        .C2(n82), .O(n539) );
  AO222CHD U105 ( .A1(N92), .A2(n79), .B1(i_round[4]), .B2(n83), .C1(N78), 
        .C2(n82), .O(n538) );
  NR2BHD U106 ( .I1(n87), .I2(n88), .O(n82) );
  INVCHD U107 ( .I(n84), .O(n83) );
  ND3CHD U108 ( .I1(n88), .I2(n86), .I3(n89), .O(n84) );
  ND2CHD U109 ( .I1(n90), .I2(n86), .O(n88) );
  OAI12CHD U110 ( .B1(n91), .B2(n92), .A1(i_round[5]), .O(n90) );
  INVCHD U111 ( .I(n89), .O(n79) );
  OAI112BHD U112 ( .C1(n93), .C2(n92), .A1(n87), .B1(n86), .O(n89) );
  INVCHD U113 ( .I(reset), .O(n86) );
  INVCHD U114 ( .I(ed), .O(n87) );
  AO12CHD U115 ( .B1(dx0[6]), .B2(n94), .A1(n95), .O(n537) );
  AO12CHD U116 ( .B1(dx0[5]), .B2(n94), .A1(n96), .O(n536) );
  AO12CHD U117 ( .B1(dx0[4]), .B2(n94), .A1(n97), .O(n535) );
  AO12CHD U118 ( .B1(dx0[3]), .B2(n94), .A1(n98), .O(n534) );
  AO12CHD U119 ( .B1(dx0[2]), .B2(n94), .A1(n99), .O(n533) );
  AO12CHD U120 ( .B1(dx0[1]), .B2(n94), .A1(n100), .O(n532) );
  OR3B2CHD U121 ( .I1(n101), .B1(n102), .B2(n103), .O(n531) );
  AOI112BHD U122 ( .C1(dx0[0]), .C2(n94), .A1(n104), .B1(n105), .O(n103) );
  INVCHD U123 ( .I(n106), .O(n105) );
  AO12CHD U124 ( .B1(dx1[6]), .B2(n94), .A1(n107), .O(n530) );
  AO12CHD U125 ( .B1(dx1[5]), .B2(n94), .A1(n95), .O(n529) );
  AO12CHD U126 ( .B1(dx1[4]), .B2(n94), .A1(n96), .O(n528) );
  AO12CHD U127 ( .B1(dx1[3]), .B2(n94), .A1(n97), .O(n527) );
  AO12CHD U128 ( .B1(dx1[2]), .B2(n94), .A1(n98), .O(n526) );
  AO12CHD U129 ( .B1(dx1[1]), .B2(n94), .A1(n99), .O(n525) );
  AO12CHD U130 ( .B1(dx1[0]), .B2(n94), .A1(n100), .O(n524) );
  OAI112BHD U131 ( .C1(n108), .C2(n109), .A1(n110), .B1(n111), .O(n100) );
  AN3B2BHD U132 ( .I1(n112), .B1(n113), .B2(n114), .O(n111) );
  NR2BHD U133 ( .I1(n115), .I2(n116), .O(n110) );
  AO12CHD U134 ( .B1(dx2[6]), .B2(n94), .A1(n117), .O(n523) );
  AO12CHD U135 ( .B1(dx2[5]), .B2(n94), .A1(n107), .O(n522) );
  AO12CHD U136 ( .B1(dx2[4]), .B2(n94), .A1(n95), .O(n521) );
  AO12CHD U137 ( .B1(dx2[3]), .B2(n94), .A1(n96), .O(n520) );
  AO12CHD U138 ( .B1(dx2[2]), .B2(n94), .A1(n97), .O(n519) );
  AO12CHD U139 ( .B1(dx2[1]), .B2(n94), .A1(n98), .O(n518) );
  AO12CHD U140 ( .B1(dx2[0]), .B2(n94), .A1(n99), .O(n517) );
  ND6EHD U141 ( .I1(n29), .I2(n118), .I3(n119), .I4(n120), .I5(n121), .I6(n122), .O(n99) );
  AOI112BHD U142 ( .C1(n123), .C2(n124), .A1(n125), .B1(n10), .O(n122) );
  OAI112BHD U143 ( .C1(n127), .C2(n128), .A1(n129), .B1(n130), .O(n125) );
  INVCHD U144 ( .I(n116), .O(n130) );
  OAI12CHD U145 ( .B1(n131), .B2(n132), .A1(n133), .O(n129) );
  ND6EHD U146 ( .I1(n119), .I2(n134), .I3(n135), .I4(n136), .I5(n13), .I6(n137), .O(n516) );
  AN4B1BHD U147 ( .I1(n106), .I2(n138), .I3(n139), .B1(n140), .O(n137) );
  AOI22BHD U148 ( .A1(dx3[6]), .A2(n94), .B1(n141), .B2(n142), .O(n139) );
  OA12CHD U149 ( .B1(n144), .B2(n145), .A1(n18), .O(n119) );
  AO12CHD U150 ( .B1(dx3[5]), .B2(n94), .A1(n117), .O(n515) );
  ND6EHD U151 ( .I1(n120), .I2(n28), .I3(n135), .I4(n24), .I5(n146), .I6(n147), 
        .O(n117) );
  AOI12CHD U152 ( .B1(n131), .B2(n142), .A1(n115), .O(n147) );
  OA112CHD U153 ( .C1(n148), .C2(n149), .A1(n150), .B1(n151), .O(n135) );
  NR2BHD U154 ( .I1(n152), .I2(n153), .O(n151) );
  AO12CHD U155 ( .B1(dx3[4]), .B2(n94), .A1(n107), .O(n514) );
  OAI112BHD U156 ( .C1(n93), .C2(n145), .A1(n53), .B1(n154), .O(n107) );
  NR2BHD U157 ( .I1(n155), .I2(n101), .O(n154) );
  OAI112BHD U158 ( .C1(n156), .C2(n144), .A1(n57), .B1(n157), .O(n101) );
  NR3BHD U159 ( .I1(n140), .I2(n158), .I3(n159), .O(n157) );
  AO12CHD U160 ( .B1(dx3[3]), .B2(n94), .A1(n95), .O(n513) );
  AO12CHD U161 ( .B1(dx3[2]), .B2(n94), .A1(n96), .O(n512) );
  ND6EHD U162 ( .I1(n35), .I2(n9), .I3(n160), .I4(n23), .I5(n112), .I6(n161), 
        .O(n96) );
  AOI112BHD U163 ( .C1(n162), .C2(n124), .A1(n163), .B1(n164), .O(n161) );
  OR3B2CHD U164 ( .I1(n159), .B1(n165), .B2(n150), .O(n163) );
  INVCHD U165 ( .I(n166), .O(n165) );
  AOI12CHD U166 ( .B1(n124), .B2(n167), .A1(n153), .O(n112) );
  AO12CHD U167 ( .B1(dx3[1]), .B2(n94), .A1(n97), .O(n511) );
  ND6EHD U168 ( .I1(n25), .I2(n160), .I3(n17), .I4(n118), .I5(n168), .I6(n169), 
        .O(n97) );
  NR2BHD U169 ( .I1(n170), .I2(n152), .O(n169) );
  AO12CHD U170 ( .B1(n109), .B2(n171), .A1(n108), .O(n168) );
  AO12CHD U171 ( .B1(dx3[0]), .B2(n94), .A1(n98), .O(n510) );
  OAI112BHD U172 ( .C1(n93), .C2(n171), .A1(n102), .B1(n172), .O(n98) );
  NR2BHD U173 ( .I1(n155), .I2(n27), .O(n172) );
  ND3CHD U174 ( .I1(n173), .I2(n174), .I3(n175), .O(n155) );
  AN3B2BHD U175 ( .I1(n138), .B1(n170), .B2(n153), .O(n175) );
  AN3B2BHD U176 ( .I1(n176), .B1(n116), .B2(n115), .O(n102) );
  NR2BHD U177 ( .I1(n36), .I2(n42), .O(n176) );
  NR3BHD U178 ( .I1(n181), .I2(n164), .I3(n140), .O(n180) );
  OAI12CHD U179 ( .B1(n149), .B2(n145), .A1(n160), .O(n181) );
  OA12CHD U180 ( .B1(n108), .B2(n145), .A1(n173), .O(n160) );
  NR2BHD U181 ( .I1(n142), .I2(n124), .O(n108) );
  AN4B1BHD U182 ( .I1(n57), .I2(n146), .I3(n134), .B1(n95), .O(n179) );
  ND2CHD U183 ( .I1(n182), .I2(n183), .O(n95) );
  AOI112BHD U184 ( .C1(n123), .C2(n184), .A1(n185), .B1(n166), .O(n183) );
  OAI22CHD U185 ( .A1(n93), .A2(n109), .B1(n128), .B2(n149), .O(n185) );
  INVCHD U186 ( .I(n162), .O(n128) );
  INVCHD U187 ( .I(n127), .O(n184) );
  NR2BHD U188 ( .I1(n186), .I2(n124), .O(n127) );
  AN4B1BHD U189 ( .I1(n32), .I2(n48), .I3(n51), .B1(n114), .O(n182) );
  ND6EHD U190 ( .I1(n118), .I2(n9), .I3(n53), .I4(n138), .I5(n187), .I6(n106), 
        .O(n114) );
  AOI12CHD U191 ( .B1(n133), .B2(n162), .A1(n116), .O(n146) );
  OR3B2CHD U192 ( .I1(n190), .B1(n191), .B2(n192), .O(n509) );
  NR3BHD U193 ( .I1(n193), .I2(n194), .I3(n195), .O(n192) );
  OAI22CHD U194 ( .A1(n20), .A2(n196), .B1(n23), .B2(n197), .O(n195) );
  OAI222BHD U195 ( .A1(n51), .A2(n198), .B1(n121), .B2(n199), .C1(n48), .C2(
        n200), .O(n194) );
  AO2222BHD U196 ( .A1(MK[95]), .A2(n27), .B1(MK[55]), .B2(n42), .C1(MK[23]), 
        .C2(n55), .D1(MK[119]), .D2(n12), .O(n193) );
  OA2222CHD U197 ( .A1(n9), .A2(n201), .B1(n118), .B2(n202), .C1(n32), .C2(
        n203), .D1(n120), .D2(n204), .O(n191) );
  AO2222BHD U198 ( .A1(mkx0[7]), .A2(n61), .B1(MK[7]), .B2(n188), .C1(MK[39]), 
        .C2(n36), .D1(MK[71]), .D2(n67), .O(n190) );
  OR3B2CHD U199 ( .I1(n207), .B1(n208), .B2(n209), .O(n508) );
  NR3BHD U200 ( .I1(n210), .I2(n211), .I3(n212), .O(n209) );
  OAI22CHD U201 ( .A1(n20), .A2(n213), .B1(n23), .B2(n214), .O(n212) );
  OAI222BHD U202 ( .A1(n51), .A2(n215), .B1(n121), .B2(n216), .C1(n48), .C2(
        n217), .O(n211) );
  AO2222BHD U203 ( .A1(MK[94]), .A2(n27), .B1(MK[54]), .B2(n42), .C1(MK[22]), 
        .C2(n56), .D1(MK[118]), .D2(n143), .O(n210) );
  OA2222CHD U204 ( .A1(n9), .A2(n218), .B1(n118), .B2(n219), .C1(n32), .C2(
        n220), .D1(n120), .D2(n221), .O(n208) );
  AO2222BHD U205 ( .A1(mkx0[6]), .A2(n61), .B1(MK[6]), .B2(n188), .C1(MK[38]), 
        .C2(n36), .D1(MK[70]), .D2(n67), .O(n207) );
  OR3B2CHD U206 ( .I1(n222), .B1(n223), .B2(n224), .O(n507) );
  NR3BHD U207 ( .I1(n225), .I2(n226), .I3(n227), .O(n224) );
  OAI22CHD U208 ( .A1(n19), .A2(n228), .B1(n23), .B2(n229), .O(n227) );
  OAI222BHD U209 ( .A1(n51), .A2(n230), .B1(n121), .B2(n231), .C1(n48), .C2(
        n232), .O(n226) );
  AO2222BHD U210 ( .A1(MK[93]), .A2(n27), .B1(MK[53]), .B2(n41), .C1(MK[21]), 
        .C2(n56), .D1(MK[117]), .D2(n12), .O(n225) );
  OA2222CHD U211 ( .A1(n9), .A2(n233), .B1(n118), .B2(n234), .C1(n32), .C2(
        n235), .D1(n120), .D2(n236), .O(n223) );
  AO2222BHD U212 ( .A1(mkx0[5]), .A2(n61), .B1(MK[5]), .B2(n52), .C1(MK[37]), 
        .C2(n36), .D1(MK[69]), .D2(n67), .O(n222) );
  OR3B2CHD U213 ( .I1(n237), .B1(n238), .B2(n239), .O(n506) );
  NR3BHD U214 ( .I1(n240), .I2(n241), .I3(n242), .O(n239) );
  OAI22CHD U215 ( .A1(n19), .A2(n243), .B1(n23), .B2(n244), .O(n242) );
  OAI222BHD U216 ( .A1(n51), .A2(n245), .B1(n121), .B2(n246), .C1(n48), .C2(
        n247), .O(n241) );
  AO2222BHD U217 ( .A1(MK[92]), .A2(n27), .B1(MK[52]), .B2(n41), .C1(MK[20]), 
        .C2(n56), .D1(MK[116]), .D2(n12), .O(n240) );
  OA2222CHD U218 ( .A1(n9), .A2(n248), .B1(n118), .B2(n249), .C1(n32), .C2(
        n250), .D1(n120), .D2(n251), .O(n238) );
  AO2222BHD U219 ( .A1(mkx0[4]), .A2(n61), .B1(MK[4]), .B2(n188), .C1(MK[36]), 
        .C2(n36), .D1(MK[68]), .D2(n67), .O(n237) );
  OR3B2CHD U220 ( .I1(n252), .B1(n253), .B2(n254), .O(n505) );
  NR3BHD U221 ( .I1(n255), .I2(n256), .I3(n257), .O(n254) );
  OAI22CHD U222 ( .A1(n19), .A2(n258), .B1(n23), .B2(n259), .O(n257) );
  OAI222BHD U223 ( .A1(n51), .A2(n260), .B1(n121), .B2(n261), .C1(n48), .C2(
        n262), .O(n256) );
  AO2222BHD U224 ( .A1(MK[91]), .A2(n27), .B1(MK[51]), .B2(n41), .C1(MK[19]), 
        .C2(n56), .D1(MK[115]), .D2(n12), .O(n255) );
  OA2222CHD U225 ( .A1(n9), .A2(n263), .B1(n118), .B2(n264), .C1(n32), .C2(
        n265), .D1(n120), .D2(n266), .O(n253) );
  AO2222BHD U226 ( .A1(mkx0[3]), .A2(n61), .B1(MK[3]), .B2(n52), .C1(MK[35]), 
        .C2(n36), .D1(MK[67]), .D2(n67), .O(n252) );
  OR3B2CHD U227 ( .I1(n267), .B1(n268), .B2(n269), .O(n504) );
  NR3BHD U228 ( .I1(n270), .I2(n271), .I3(n272), .O(n269) );
  OAI22CHD U229 ( .A1(n19), .A2(n273), .B1(n24), .B2(n274), .O(n272) );
  OAI222BHD U230 ( .A1(n51), .A2(n275), .B1(n121), .B2(n276), .C1(n48), .C2(
        n277), .O(n271) );
  AO2222BHD U231 ( .A1(MK[90]), .A2(n27), .B1(MK[50]), .B2(n41), .C1(MK[18]), 
        .C2(n56), .D1(MK[114]), .D2(n12), .O(n270) );
  OA2222CHD U232 ( .A1(n9), .A2(n278), .B1(n118), .B2(n279), .C1(n32), .C2(
        n280), .D1(n120), .D2(n281), .O(n268) );
  AO2222BHD U233 ( .A1(mkx0[2]), .A2(n61), .B1(MK[2]), .B2(n188), .C1(MK[34]), 
        .C2(n36), .D1(MK[66]), .D2(n67), .O(n267) );
  OR3B2CHD U234 ( .I1(n282), .B1(n283), .B2(n284), .O(n503) );
  NR3BHD U235 ( .I1(n285), .I2(n286), .I3(n287), .O(n284) );
  OAI22CHD U236 ( .A1(n19), .A2(n288), .B1(n23), .B2(n289), .O(n287) );
  OAI222BHD U237 ( .A1(n51), .A2(n290), .B1(n121), .B2(n291), .C1(n48), .C2(
        n292), .O(n286) );
  AO2222BHD U238 ( .A1(MK[89]), .A2(n27), .B1(MK[49]), .B2(n41), .C1(MK[17]), 
        .C2(n56), .D1(MK[113]), .D2(n12), .O(n285) );
  OA2222CHD U239 ( .A1(n9), .A2(n293), .B1(n118), .B2(n294), .C1(n33), .C2(
        n295), .D1(n120), .D2(n296), .O(n283) );
  AO2222BHD U240 ( .A1(mkx0[1]), .A2(n61), .B1(MK[1]), .B2(n188), .C1(MK[33]), 
        .C2(n36), .D1(MK[65]), .D2(n67), .O(n282) );
  OR3B2CHD U241 ( .I1(n297), .B1(n298), .B2(n299), .O(n502) );
  NR3BHD U242 ( .I1(n300), .I2(n301), .I3(n302), .O(n299) );
  OAI22CHD U243 ( .A1(n19), .A2(n303), .B1(n23), .B2(n304), .O(n302) );
  OAI222BHD U244 ( .A1(n51), .A2(n305), .B1(n121), .B2(n306), .C1(n48), .C2(
        n307), .O(n301) );
  AO2222BHD U245 ( .A1(MK[88]), .A2(n27), .B1(MK[48]), .B2(n41), .C1(MK[16]), 
        .C2(n56), .D1(MK[112]), .D2(n12), .O(n300) );
  OA2222CHD U246 ( .A1(n9), .A2(n308), .B1(n118), .B2(n309), .C1(n32), .C2(
        n310), .D1(n120), .D2(n311), .O(n298) );
  AO2222BHD U247 ( .A1(mkx0[0]), .A2(n61), .B1(MK[0]), .B2(n188), .C1(MK[32]), 
        .C2(n36), .D1(MK[64]), .D2(n67), .O(n297) );
  OR3B2CHD U248 ( .I1(n312), .B1(n313), .B2(n314), .O(n501) );
  NR3BHD U249 ( .I1(n315), .I2(n316), .I3(n317), .O(n314) );
  OAI22CHD U250 ( .A1(n19), .A2(n318), .B1(n23), .B2(n198), .O(n317) );
  OAI222BHD U251 ( .A1(n51), .A2(n319), .B1(n121), .B2(n320), .C1(n48), .C2(
        n321), .O(n316) );
  AO2222BHD U252 ( .A1(MK[103]), .A2(n27), .B1(MK[63]), .B2(n41), .C1(MK[31]), 
        .C2(n56), .D1(MK[127]), .D2(n12), .O(n315) );
  OA2222CHD U253 ( .A1(n9), .A2(n196), .B1(n118), .B2(n322), .C1(n32), .C2(
        n323), .D1(n120), .D2(n324), .O(n313) );
  AO2222BHD U254 ( .A1(mkx1[7]), .A2(n61), .B1(MK[15]), .B2(n188), .C1(MK[47]), 
        .C2(n36), .D1(MK[79]), .D2(n67), .O(n312) );
  OR3B2CHD U255 ( .I1(n325), .B1(n326), .B2(n327), .O(n500) );
  NR3BHD U256 ( .I1(n328), .I2(n329), .I3(n330), .O(n327) );
  OAI22CHD U257 ( .A1(n19), .A2(n331), .B1(n23), .B2(n215), .O(n330) );
  OAI222BHD U258 ( .A1(n51), .A2(n332), .B1(n121), .B2(n333), .C1(n48), .C2(
        n334), .O(n329) );
  AO2222BHD U259 ( .A1(MK[102]), .A2(n27), .B1(MK[62]), .B2(n41), .C1(MK[30]), 
        .C2(n56), .D1(MK[126]), .D2(n12), .O(n328) );
  OA2222CHD U260 ( .A1(n126), .A2(n213), .B1(n118), .B2(n335), .C1(n32), .C2(
        n336), .D1(n120), .D2(n337), .O(n326) );
  AO2222BHD U261 ( .A1(mkx1[6]), .A2(n61), .B1(MK[14]), .B2(n188), .C1(MK[46]), 
        .C2(n36), .D1(MK[78]), .D2(n67), .O(n325) );
  OR3B2CHD U262 ( .I1(n338), .B1(n339), .B2(n340), .O(n499) );
  NR3BHD U263 ( .I1(n341), .I2(n342), .I3(n343), .O(n340) );
  OAI22CHD U264 ( .A1(n19), .A2(n344), .B1(n24), .B2(n230), .O(n343) );
  OAI222BHD U265 ( .A1(n50), .A2(n345), .B1(n121), .B2(n346), .C1(n47), .C2(
        n347), .O(n342) );
  AO2222BHD U266 ( .A1(MK[101]), .A2(n27), .B1(MK[61]), .B2(n41), .C1(MK[29]), 
        .C2(n56), .D1(MK[125]), .D2(n12), .O(n341) );
  OA2222CHD U267 ( .A1(n126), .A2(n228), .B1(n118), .B2(n348), .C1(n33), .C2(
        n349), .D1(n120), .D2(n350), .O(n339) );
  AO2222BHD U268 ( .A1(mkx1[5]), .A2(n62), .B1(MK[13]), .B2(n188), .C1(MK[45]), 
        .C2(n37), .D1(MK[77]), .D2(n68), .O(n338) );
  OR3B2CHD U269 ( .I1(n351), .B1(n352), .B2(n353), .O(n498) );
  NR3BHD U270 ( .I1(n354), .I2(n355), .I3(n356), .O(n353) );
  OAI22CHD U271 ( .A1(n19), .A2(n357), .B1(n24), .B2(n245), .O(n356) );
  OAI222BHD U272 ( .A1(n50), .A2(n358), .B1(n121), .B2(n359), .C1(n47), .C2(
        n360), .O(n355) );
  AO2222BHD U273 ( .A1(MK[100]), .A2(n27), .B1(MK[60]), .B2(n41), .C1(MK[28]), 
        .C2(n56), .D1(MK[124]), .D2(n12), .O(n354) );
  OA2222CHD U274 ( .A1(n126), .A2(n243), .B1(n118), .B2(n361), .C1(n33), .C2(
        n362), .D1(n120), .D2(n363), .O(n352) );
  AO2222BHD U275 ( .A1(mkx1[4]), .A2(n62), .B1(MK[12]), .B2(n188), .C1(MK[44]), 
        .C2(n37), .D1(MK[76]), .D2(n68), .O(n351) );
  OR3B2CHD U276 ( .I1(n364), .B1(n365), .B2(n366), .O(n497) );
  NR3BHD U277 ( .I1(n367), .I2(n368), .I3(n369), .O(n366) );
  OAI22CHD U278 ( .A1(n18), .A2(n370), .B1(n24), .B2(n260), .O(n369) );
  OAI222BHD U279 ( .A1(n50), .A2(n371), .B1(n121), .B2(n372), .C1(n47), .C2(
        n373), .O(n368) );
  AO2222BHD U280 ( .A1(MK[99]), .A2(n27), .B1(MK[59]), .B2(n40), .C1(MK[27]), 
        .C2(n55), .D1(MK[123]), .D2(n12), .O(n367) );
  OA2222CHD U281 ( .A1(n126), .A2(n258), .B1(n118), .B2(n374), .C1(n33), .C2(
        n375), .D1(n120), .D2(n376), .O(n365) );
  AO2222BHD U282 ( .A1(mkx1[3]), .A2(n62), .B1(MK[11]), .B2(n188), .C1(MK[43]), 
        .C2(n37), .D1(MK[75]), .D2(n68), .O(n364) );
  OR3B2CHD U283 ( .I1(n377), .B1(n378), .B2(n379), .O(n496) );
  NR3BHD U284 ( .I1(n380), .I2(n381), .I3(n382), .O(n379) );
  OAI22CHD U285 ( .A1(n18), .A2(n383), .B1(n24), .B2(n275), .O(n382) );
  OAI222BHD U286 ( .A1(n50), .A2(n384), .B1(n121), .B2(n385), .C1(n47), .C2(
        n386), .O(n381) );
  AO2222BHD U287 ( .A1(MK[98]), .A2(n27), .B1(MK[58]), .B2(n40), .C1(MK[26]), 
        .C2(n55), .D1(MK[122]), .D2(n12), .O(n380) );
  OA2222CHD U288 ( .A1(n126), .A2(n273), .B1(n118), .B2(n387), .C1(n33), .C2(
        n388), .D1(n120), .D2(n389), .O(n378) );
  AO2222BHD U289 ( .A1(mkx1[2]), .A2(n62), .B1(MK[10]), .B2(n188), .C1(MK[42]), 
        .C2(n37), .D1(MK[74]), .D2(n68), .O(n377) );
  OR3B2CHD U290 ( .I1(n390), .B1(n391), .B2(n392), .O(n495) );
  NR3BHD U291 ( .I1(n393), .I2(n394), .I3(n395), .O(n392) );
  OAI22CHD U292 ( .A1(n18), .A2(n396), .B1(n24), .B2(n290), .O(n395) );
  OAI222BHD U293 ( .A1(n50), .A2(n397), .B1(n121), .B2(n398), .C1(n47), .C2(
        n399), .O(n394) );
  AO2222BHD U294 ( .A1(MK[97]), .A2(n27), .B1(MK[57]), .B2(n40), .C1(MK[25]), 
        .C2(n55), .D1(MK[121]), .D2(n12), .O(n393) );
  OA2222CHD U295 ( .A1(n126), .A2(n288), .B1(n118), .B2(n400), .C1(n33), .C2(
        n401), .D1(n120), .D2(n402), .O(n391) );
  AO2222BHD U296 ( .A1(mkx1[1]), .A2(n62), .B1(MK[9]), .B2(n188), .C1(MK[41]), 
        .C2(n37), .D1(MK[73]), .D2(n68), .O(n390) );
  OR3B2CHD U297 ( .I1(n403), .B1(n404), .B2(n405), .O(n494) );
  NR3BHD U298 ( .I1(n406), .I2(n407), .I3(n408), .O(n405) );
  OAI22CHD U299 ( .A1(n18), .A2(n409), .B1(n24), .B2(n305), .O(n408) );
  OAI222BHD U300 ( .A1(n50), .A2(n410), .B1(n121), .B2(n411), .C1(n47), .C2(
        n412), .O(n407) );
  AO2222BHD U301 ( .A1(MK[96]), .A2(n27), .B1(MK[56]), .B2(n40), .C1(MK[24]), 
        .C2(n55), .D1(MK[120]), .D2(n143), .O(n406) );
  OA2222CHD U302 ( .A1(n126), .A2(n303), .B1(n118), .B2(n413), .C1(n33), .C2(
        n414), .D1(n120), .D2(n415), .O(n404) );
  AO2222BHD U303 ( .A1(mkx1[0]), .A2(n62), .B1(MK[8]), .B2(n188), .C1(MK[40]), 
        .C2(n37), .D1(MK[72]), .D2(n68), .O(n403) );
  OR3B2CHD U304 ( .I1(n416), .B1(n417), .B2(n418), .O(n493) );
  NR3BHD U305 ( .I1(n419), .I2(n420), .I3(n421), .O(n418) );
  OAI22CHD U306 ( .A1(n18), .A2(n204), .B1(n24), .B2(n319), .O(n421) );
  INVCHD U307 ( .I(MK[95]), .O(n319) );
  OAI222BHD U308 ( .A1(n50), .A2(n201), .B1(n121), .B2(n202), .C1(n47), .C2(
        n203), .O(n420) );
  INVCHD U309 ( .I(MK[31]), .O(n203) );
  INVCHD U310 ( .I(MK[63]), .O(n202) );
  AO2222BHD U311 ( .A1(MK[111]), .A2(n27), .B1(MK[7]), .B2(n40), .C1(MK[39]), 
        .C2(n55), .D1(MK[71]), .D2(n143), .O(n419) );
  OA2222CHD U312 ( .A1(n126), .A2(n318), .B1(n118), .B2(n200), .C1(n33), .C2(
        n199), .D1(n120), .D2(n197), .O(n417) );
  INVCHD U313 ( .I(MK[79]), .O(n197) );
  INVCHD U314 ( .I(MK[47]), .O(n199) );
  INVCHD U315 ( .I(MK[15]), .O(n200) );
  INVCHD U316 ( .I(MK[119]), .O(n318) );
  AO2222BHD U317 ( .A1(mkx2[7]), .A2(n62), .B1(MK[23]), .B2(n188), .C1(MK[55]), 
        .C2(n37), .D1(MK[87]), .D2(n68), .O(n416) );
  OR3B2CHD U318 ( .I1(n422), .B1(n423), .B2(n424), .O(n492) );
  NR3BHD U319 ( .I1(n425), .I2(n426), .I3(n427), .O(n424) );
  OAI22CHD U320 ( .A1(n18), .A2(n221), .B1(n24), .B2(n332), .O(n427) );
  INVCHD U321 ( .I(MK[94]), .O(n332) );
  OAI222BHD U322 ( .A1(n50), .A2(n218), .B1(n121), .B2(n219), .C1(n47), .C2(
        n220), .O(n426) );
  INVCHD U323 ( .I(MK[30]), .O(n220) );
  INVCHD U324 ( .I(MK[62]), .O(n219) );
  AO2222BHD U325 ( .A1(MK[110]), .A2(n27), .B1(MK[6]), .B2(n40), .C1(MK[38]), 
        .C2(n55), .D1(MK[70]), .D2(n143), .O(n425) );
  OA2222CHD U326 ( .A1(n126), .A2(n331), .B1(n118), .B2(n217), .C1(n33), .C2(
        n216), .D1(n120), .D2(n214), .O(n423) );
  INVCHD U327 ( .I(MK[78]), .O(n214) );
  INVCHD U328 ( .I(MK[46]), .O(n216) );
  INVCHD U329 ( .I(MK[14]), .O(n217) );
  INVCHD U330 ( .I(MK[118]), .O(n331) );
  AO2222BHD U331 ( .A1(mkx2[6]), .A2(n62), .B1(MK[22]), .B2(n188), .C1(MK[54]), 
        .C2(n37), .D1(MK[86]), .D2(n68), .O(n422) );
  OR3B2CHD U332 ( .I1(n428), .B1(n429), .B2(n430), .O(n491) );
  NR3BHD U333 ( .I1(n431), .I2(n432), .I3(n433), .O(n430) );
  OAI22CHD U334 ( .A1(n18), .A2(n236), .B1(n24), .B2(n345), .O(n433) );
  INVCHD U335 ( .I(MK[93]), .O(n345) );
  OAI222BHD U336 ( .A1(n50), .A2(n233), .B1(n121), .B2(n234), .C1(n47), .C2(
        n235), .O(n432) );
  INVCHD U337 ( .I(MK[29]), .O(n235) );
  INVCHD U338 ( .I(MK[61]), .O(n234) );
  AO2222BHD U339 ( .A1(MK[109]), .A2(n27), .B1(MK[5]), .B2(n40), .C1(MK[37]), 
        .C2(n55), .D1(MK[69]), .D2(n143), .O(n431) );
  OA2222CHD U340 ( .A1(n126), .A2(n344), .B1(n118), .B2(n232), .C1(n33), .C2(
        n231), .D1(n120), .D2(n229), .O(n429) );
  INVCHD U341 ( .I(MK[77]), .O(n229) );
  INVCHD U342 ( .I(MK[45]), .O(n231) );
  INVCHD U343 ( .I(MK[13]), .O(n232) );
  INVCHD U344 ( .I(MK[117]), .O(n344) );
  AO2222BHD U345 ( .A1(mkx2[5]), .A2(n62), .B1(MK[21]), .B2(n188), .C1(MK[53]), 
        .C2(n37), .D1(MK[85]), .D2(n68), .O(n428) );
  OR3B2CHD U346 ( .I1(n434), .B1(n435), .B2(n436), .O(n490) );
  NR3BHD U347 ( .I1(n437), .I2(n438), .I3(n439), .O(n436) );
  OAI22CHD U348 ( .A1(n18), .A2(n251), .B1(n25), .B2(n358), .O(n439) );
  INVCHD U349 ( .I(MK[92]), .O(n358) );
  OAI222BHD U350 ( .A1(n50), .A2(n248), .B1(n121), .B2(n249), .C1(n47), .C2(
        n250), .O(n438) );
  INVCHD U351 ( .I(MK[28]), .O(n250) );
  INVCHD U352 ( .I(MK[60]), .O(n249) );
  AO2222BHD U353 ( .A1(MK[108]), .A2(n27), .B1(MK[4]), .B2(n40), .C1(MK[36]), 
        .C2(n55), .D1(MK[68]), .D2(n143), .O(n437) );
  OA2222CHD U354 ( .A1(n126), .A2(n357), .B1(n118), .B2(n247), .C1(n34), .C2(
        n246), .D1(n120), .D2(n244), .O(n435) );
  INVCHD U355 ( .I(MK[76]), .O(n244) );
  INVCHD U356 ( .I(MK[44]), .O(n246) );
  INVCHD U357 ( .I(MK[12]), .O(n247) );
  INVCHD U358 ( .I(MK[116]), .O(n357) );
  AO2222BHD U359 ( .A1(mkx2[4]), .A2(n62), .B1(MK[20]), .B2(n188), .C1(MK[52]), 
        .C2(n37), .D1(MK[84]), .D2(n68), .O(n434) );
  OR3B2CHD U360 ( .I1(n440), .B1(n441), .B2(n442), .O(n489) );
  NR3BHD U361 ( .I1(n443), .I2(n444), .I3(n445), .O(n442) );
  OAI22CHD U362 ( .A1(n18), .A2(n266), .B1(n25), .B2(n371), .O(n445) );
  INVCHD U363 ( .I(MK[91]), .O(n371) );
  OAI222BHD U364 ( .A1(n50), .A2(n263), .B1(n121), .B2(n264), .C1(n47), .C2(
        n265), .O(n444) );
  INVCHD U365 ( .I(MK[27]), .O(n265) );
  INVCHD U366 ( .I(MK[59]), .O(n264) );
  AO2222BHD U367 ( .A1(MK[107]), .A2(n27), .B1(MK[3]), .B2(n40), .C1(MK[35]), 
        .C2(n55), .D1(MK[67]), .D2(n143), .O(n443) );
  OA2222CHD U368 ( .A1(n126), .A2(n370), .B1(n118), .B2(n262), .C1(n34), .C2(
        n261), .D1(n120), .D2(n259), .O(n441) );
  INVCHD U369 ( .I(MK[75]), .O(n259) );
  INVCHD U370 ( .I(MK[43]), .O(n261) );
  INVCHD U371 ( .I(MK[11]), .O(n262) );
  INVCHD U372 ( .I(MK[115]), .O(n370) );
  AO2222BHD U373 ( .A1(mkx2[3]), .A2(n63), .B1(MK[19]), .B2(n188), .C1(MK[51]), 
        .C2(n37), .D1(MK[83]), .D2(n69), .O(n440) );
  OR3B2CHD U374 ( .I1(n446), .B1(n447), .B2(n448), .O(n488) );
  NR3BHD U375 ( .I1(n449), .I2(n450), .I3(n451), .O(n448) );
  OAI22CHD U376 ( .A1(n18), .A2(n281), .B1(n25), .B2(n384), .O(n451) );
  INVCHD U377 ( .I(MK[90]), .O(n384) );
  OAI222BHD U378 ( .A1(n49), .A2(n278), .B1(n121), .B2(n279), .C1(n46), .C2(
        n280), .O(n450) );
  INVCHD U379 ( .I(MK[26]), .O(n280) );
  INVCHD U380 ( .I(MK[58]), .O(n279) );
  AO2222BHD U381 ( .A1(MK[106]), .A2(n27), .B1(MK[2]), .B2(n40), .C1(MK[34]), 
        .C2(n55), .D1(MK[66]), .D2(n143), .O(n449) );
  OA2222CHD U382 ( .A1(n126), .A2(n383), .B1(n118), .B2(n277), .C1(n34), .C2(
        n276), .D1(n120), .D2(n274), .O(n447) );
  INVCHD U383 ( .I(MK[74]), .O(n274) );
  INVCHD U384 ( .I(MK[42]), .O(n276) );
  INVCHD U385 ( .I(MK[10]), .O(n277) );
  INVCHD U386 ( .I(MK[114]), .O(n383) );
  AO2222BHD U387 ( .A1(mkx2[2]), .A2(n63), .B1(MK[18]), .B2(n188), .C1(MK[50]), 
        .C2(n38), .D1(MK[82]), .D2(n69), .O(n446) );
  OR3B2CHD U388 ( .I1(n452), .B1(n453), .B2(n454), .O(n487) );
  NR3BHD U389 ( .I1(n455), .I2(n456), .I3(n457), .O(n454) );
  OAI22CHD U390 ( .A1(n17), .A2(n296), .B1(n25), .B2(n397), .O(n457) );
  INVCHD U391 ( .I(MK[89]), .O(n397) );
  OAI222BHD U392 ( .A1(n49), .A2(n293), .B1(n121), .B2(n294), .C1(n46), .C2(
        n295), .O(n456) );
  INVCHD U393 ( .I(MK[25]), .O(n295) );
  INVCHD U394 ( .I(MK[57]), .O(n294) );
  AO2222BHD U395 ( .A1(MK[105]), .A2(n27), .B1(MK[1]), .B2(n39), .C1(MK[33]), 
        .C2(n55), .D1(MK[65]), .D2(n12), .O(n455) );
  OA2222CHD U396 ( .A1(n126), .A2(n396), .B1(n118), .B2(n292), .C1(n34), .C2(
        n291), .D1(n120), .D2(n289), .O(n453) );
  INVCHD U397 ( .I(MK[73]), .O(n289) );
  INVCHD U398 ( .I(MK[41]), .O(n291) );
  INVCHD U399 ( .I(MK[9]), .O(n292) );
  INVCHD U400 ( .I(MK[113]), .O(n396) );
  AO2222BHD U401 ( .A1(mkx2[1]), .A2(n63), .B1(MK[17]), .B2(n188), .C1(MK[49]), 
        .C2(n38), .D1(MK[81]), .D2(n69), .O(n452) );
  OR3B2CHD U402 ( .I1(n458), .B1(n459), .B2(n460), .O(n486) );
  NR3BHD U403 ( .I1(n461), .I2(n462), .I3(n463), .O(n460) );
  OAI22CHD U404 ( .A1(n17), .A2(n311), .B1(n25), .B2(n410), .O(n463) );
  INVCHD U405 ( .I(MK[88]), .O(n410) );
  OAI222BHD U406 ( .A1(n49), .A2(n308), .B1(n121), .B2(n309), .C1(n46), .C2(
        n310), .O(n462) );
  INVCHD U407 ( .I(MK[24]), .O(n310) );
  INVCHD U408 ( .I(MK[56]), .O(n309) );
  AO2222BHD U409 ( .A1(MK[104]), .A2(n27), .B1(MK[0]), .B2(n39), .C1(MK[32]), 
        .C2(n56), .D1(MK[64]), .D2(n12), .O(n461) );
  OA2222CHD U410 ( .A1(n126), .A2(n409), .B1(n118), .B2(n307), .C1(n34), .C2(
        n306), .D1(n120), .D2(n304), .O(n459) );
  INVCHD U411 ( .I(MK[72]), .O(n304) );
  INVCHD U412 ( .I(MK[40]), .O(n306) );
  INVCHD U413 ( .I(MK[8]), .O(n307) );
  INVCHD U414 ( .I(MK[112]), .O(n409) );
  AO2222BHD U415 ( .A1(mkx2[0]), .A2(n63), .B1(MK[16]), .B2(n188), .C1(MK[48]), 
        .C2(n38), .D1(MK[80]), .D2(n69), .O(n458) );
  OR3B2CHD U416 ( .I1(n464), .B1(n465), .B2(n466), .O(n485) );
  NR3BHD U417 ( .I1(n467), .I2(n468), .I3(n469), .O(n466) );
  OAI22CHD U418 ( .A1(n17), .A2(n324), .B1(n25), .B2(n201), .O(n469) );
  INVCHD U419 ( .I(MK[103]), .O(n201) );
  INVCHD U420 ( .I(MK[71]), .O(n324) );
  OAI222BHD U421 ( .A1(n49), .A2(n196), .B1(n121), .B2(n322), .C1(n46), .C2(
        n323), .O(n468) );
  INVCHD U422 ( .I(MK[39]), .O(n323) );
  INVCHD U423 ( .I(MK[7]), .O(n322) );
  INVCHD U424 ( .I(MK[111]), .O(n196) );
  AO2222BHD U425 ( .A1(MK[119]), .A2(n27), .B1(MK[15]), .B2(n39), .C1(MK[47]), 
        .C2(n55), .D1(MK[79]), .D2(n143), .O(n467) );
  OA2222CHD U426 ( .A1(n126), .A2(n204), .B1(n118), .B2(n321), .C1(n34), .C2(
        n320), .D1(n120), .D2(n198), .O(n465) );
  INVCHD U427 ( .I(MK[87]), .O(n198) );
  INVCHD U428 ( .I(MK[55]), .O(n320) );
  INVCHD U429 ( .I(MK[23]), .O(n321) );
  INVCHD U430 ( .I(MK[127]), .O(n204) );
  AO2222BHD U431 ( .A1(mkx3[7]), .A2(n63), .B1(MK[31]), .B2(n188), .C1(MK[63]), 
        .C2(n38), .D1(MK[95]), .D2(n69), .O(n464) );
  OR3B2CHD U432 ( .I1(n470), .B1(n471), .B2(n472), .O(n484) );
  NR3BHD U433 ( .I1(n473), .I2(n474), .I3(n475), .O(n472) );
  OAI22CHD U434 ( .A1(n17), .A2(n337), .B1(n25), .B2(n218), .O(n475) );
  INVCHD U435 ( .I(MK[102]), .O(n218) );
  INVCHD U436 ( .I(MK[70]), .O(n337) );
  OAI222BHD U437 ( .A1(n49), .A2(n213), .B1(n121), .B2(n335), .C1(n46), .C2(
        n336), .O(n474) );
  INVCHD U438 ( .I(MK[38]), .O(n336) );
  INVCHD U439 ( .I(MK[6]), .O(n335) );
  INVCHD U440 ( .I(MK[110]), .O(n213) );
  AO2222BHD U441 ( .A1(MK[118]), .A2(n27), .B1(MK[14]), .B2(n39), .C1(MK[46]), 
        .C2(n56), .D1(MK[78]), .D2(n143), .O(n473) );
  OA2222CHD U442 ( .A1(n126), .A2(n221), .B1(n118), .B2(n334), .C1(n34), .C2(
        n333), .D1(n120), .D2(n215), .O(n471) );
  INVCHD U443 ( .I(MK[86]), .O(n215) );
  INVCHD U444 ( .I(MK[54]), .O(n333) );
  INVCHD U445 ( .I(MK[22]), .O(n334) );
  INVCHD U446 ( .I(MK[126]), .O(n221) );
  AO2222BHD U447 ( .A1(mkx3[6]), .A2(n63), .B1(MK[30]), .B2(n188), .C1(MK[62]), 
        .C2(n38), .D1(MK[94]), .D2(n69), .O(n470) );
  OR3B2CHD U448 ( .I1(n476), .B1(n477), .B2(n544), .O(n483) );
  NR3BHD U449 ( .I1(n545), .I2(n546), .I3(n547), .O(n544) );
  OAI22CHD U450 ( .A1(n17), .A2(n350), .B1(n25), .B2(n233), .O(n547) );
  INVCHD U451 ( .I(MK[101]), .O(n233) );
  INVCHD U452 ( .I(MK[69]), .O(n350) );
  OAI222BHD U453 ( .A1(n49), .A2(n228), .B1(n121), .B2(n348), .C1(n46), .C2(
        n349), .O(n546) );
  INVCHD U454 ( .I(MK[37]), .O(n349) );
  INVCHD U455 ( .I(MK[5]), .O(n348) );
  INVCHD U456 ( .I(MK[109]), .O(n228) );
  AO2222BHD U457 ( .A1(MK[117]), .A2(n27), .B1(MK[13]), .B2(n39), .C1(MK[45]), 
        .C2(n55), .D1(MK[77]), .D2(n143), .O(n545) );
  OA2222CHD U458 ( .A1(n126), .A2(n236), .B1(n118), .B2(n347), .C1(n34), .C2(
        n346), .D1(n120), .D2(n230), .O(n477) );
  INVCHD U459 ( .I(MK[85]), .O(n230) );
  INVCHD U460 ( .I(MK[53]), .O(n346) );
  INVCHD U461 ( .I(MK[21]), .O(n347) );
  INVCHD U462 ( .I(MK[125]), .O(n236) );
  AO2222BHD U463 ( .A1(mkx3[5]), .A2(n63), .B1(MK[29]), .B2(n188), .C1(MK[61]), 
        .C2(n38), .D1(MK[93]), .D2(n69), .O(n476) );
  OR3B2CHD U464 ( .I1(n548), .B1(n549), .B2(n550), .O(n482) );
  NR3BHD U465 ( .I1(n551), .I2(n552), .I3(n553), .O(n550) );
  OAI22CHD U466 ( .A1(n17), .A2(n363), .B1(n25), .B2(n248), .O(n553) );
  INVCHD U467 ( .I(MK[100]), .O(n248) );
  INVCHD U468 ( .I(MK[68]), .O(n363) );
  OAI222BHD U469 ( .A1(n49), .A2(n243), .B1(n121), .B2(n361), .C1(n46), .C2(
        n362), .O(n552) );
  INVCHD U470 ( .I(MK[36]), .O(n362) );
  INVCHD U471 ( .I(MK[4]), .O(n361) );
  INVCHD U472 ( .I(MK[108]), .O(n243) );
  AO2222BHD U473 ( .A1(MK[116]), .A2(n27), .B1(MK[12]), .B2(n39), .C1(MK[44]), 
        .C2(n56), .D1(MK[76]), .D2(n143), .O(n551) );
  OA2222CHD U474 ( .A1(n126), .A2(n251), .B1(n118), .B2(n360), .C1(n34), .C2(
        n359), .D1(n120), .D2(n245), .O(n549) );
  INVCHD U475 ( .I(MK[84]), .O(n245) );
  INVCHD U476 ( .I(MK[52]), .O(n359) );
  INVCHD U477 ( .I(MK[20]), .O(n360) );
  INVCHD U478 ( .I(MK[124]), .O(n251) );
  AO2222BHD U479 ( .A1(mkx3[4]), .A2(n63), .B1(MK[28]), .B2(n188), .C1(MK[60]), 
        .C2(n38), .D1(MK[92]), .D2(n69), .O(n548) );
  OR3B2CHD U480 ( .I1(n554), .B1(n555), .B2(n556), .O(n481) );
  NR3BHD U481 ( .I1(n557), .I2(n558), .I3(n559), .O(n556) );
  OAI22CHD U482 ( .A1(n17), .A2(n376), .B1(n26), .B2(n263), .O(n559) );
  INVCHD U483 ( .I(MK[99]), .O(n263) );
  INVCHD U484 ( .I(MK[67]), .O(n376) );
  OAI222BHD U485 ( .A1(n49), .A2(n258), .B1(n121), .B2(n374), .C1(n46), .C2(
        n375), .O(n558) );
  INVCHD U486 ( .I(MK[35]), .O(n375) );
  INVCHD U487 ( .I(MK[3]), .O(n374) );
  INVCHD U488 ( .I(MK[107]), .O(n258) );
  AO2222BHD U489 ( .A1(MK[115]), .A2(n27), .B1(MK[11]), .B2(n39), .C1(MK[43]), 
        .C2(n55), .D1(MK[75]), .D2(n143), .O(n557) );
  OA2222CHD U490 ( .A1(n126), .A2(n266), .B1(n118), .B2(n373), .C1(n34), .C2(
        n372), .D1(n120), .D2(n260), .O(n555) );
  INVCHD U491 ( .I(MK[83]), .O(n260) );
  INVCHD U492 ( .I(MK[51]), .O(n372) );
  INVCHD U493 ( .I(MK[19]), .O(n373) );
  INVCHD U494 ( .I(MK[123]), .O(n266) );
  AO2222BHD U495 ( .A1(mkx3[3]), .A2(n63), .B1(MK[27]), .B2(n188), .C1(MK[59]), 
        .C2(n38), .D1(MK[91]), .D2(n69), .O(n554) );
  OR3B2CHD U496 ( .I1(n560), .B1(n561), .B2(n562), .O(n480) );
  NR3BHD U497 ( .I1(n563), .I2(n564), .I3(n565), .O(n562) );
  OAI22CHD U498 ( .A1(n17), .A2(n389), .B1(n26), .B2(n278), .O(n565) );
  INVCHD U499 ( .I(MK[98]), .O(n278) );
  INVCHD U500 ( .I(MK[66]), .O(n389) );
  OAI222BHD U501 ( .A1(n49), .A2(n273), .B1(n121), .B2(n387), .C1(n46), .C2(
        n388), .O(n564) );
  INVCHD U502 ( .I(MK[34]), .O(n388) );
  INVCHD U503 ( .I(MK[2]), .O(n387) );
  INVCHD U504 ( .I(MK[106]), .O(n273) );
  AO2222BHD U505 ( .A1(MK[114]), .A2(n27), .B1(MK[10]), .B2(n39), .C1(MK[42]), 
        .C2(n56), .D1(MK[74]), .D2(n143), .O(n563) );
  OA2222CHD U506 ( .A1(n126), .A2(n281), .B1(n118), .B2(n386), .C1(n35), .C2(
        n385), .D1(n120), .D2(n275), .O(n561) );
  INVCHD U507 ( .I(MK[82]), .O(n275) );
  INVCHD U508 ( .I(MK[50]), .O(n385) );
  INVCHD U509 ( .I(MK[18]), .O(n386) );
  INVCHD U510 ( .I(MK[122]), .O(n281) );
  AO2222BHD U511 ( .A1(mkx3[2]), .A2(n63), .B1(MK[26]), .B2(n188), .C1(MK[58]), 
        .C2(n38), .D1(MK[90]), .D2(n69), .O(n560) );
  OR3B2CHD U512 ( .I1(n566), .B1(n567), .B2(n568), .O(n479) );
  NR3BHD U513 ( .I1(n569), .I2(n570), .I3(n571), .O(n568) );
  OAI22CHD U514 ( .A1(n17), .A2(n402), .B1(n25), .B2(n293), .O(n571) );
  INVCHD U515 ( .I(MK[97]), .O(n293) );
  INVCHD U516 ( .I(MK[65]), .O(n402) );
  OAI222BHD U517 ( .A1(n49), .A2(n288), .B1(n121), .B2(n400), .C1(n46), .C2(
        n401), .O(n570) );
  INVCHD U518 ( .I(MK[33]), .O(n401) );
  INVCHD U519 ( .I(MK[1]), .O(n400) );
  INVCHD U520 ( .I(MK[105]), .O(n288) );
  AO2222BHD U521 ( .A1(MK[113]), .A2(n27), .B1(MK[9]), .B2(n39), .C1(MK[41]), 
        .C2(n55), .D1(MK[73]), .D2(n143), .O(n569) );
  OA2222CHD U522 ( .A1(n126), .A2(n296), .B1(n118), .B2(n399), .C1(n35), .C2(
        n398), .D1(n120), .D2(n290), .O(n567) );
  INVCHD U523 ( .I(MK[81]), .O(n290) );
  INVCHD U524 ( .I(MK[49]), .O(n398) );
  INVCHD U525 ( .I(MK[17]), .O(n399) );
  INVCHD U526 ( .I(MK[121]), .O(n296) );
  AO2222BHD U527 ( .A1(mkx3[1]), .A2(n64), .B1(MK[25]), .B2(n188), .C1(MK[57]), 
        .C2(n38), .D1(MK[89]), .D2(n70), .O(n566) );
  OR3B2CHD U528 ( .I1(n572), .B1(n573), .B2(n574), .O(n478) );
  NR3BHD U529 ( .I1(n575), .I2(n576), .I3(n577), .O(n574) );
  OAI22CHD U530 ( .A1(n17), .A2(n415), .B1(n23), .B2(n308), .O(n577) );
  INVCHD U531 ( .I(MK[96]), .O(n308) );
  NR2BHD U532 ( .I1(n578), .I2(n92), .O(n140) );
  INVCHD U533 ( .I(MK[64]), .O(n415) );
  INVCHD U534 ( .I(n187), .O(n158) );
  OAI222BHD U535 ( .A1(n49), .A2(n303), .B1(n121), .B2(n413), .C1(n46), .C2(
        n414), .O(n576) );
  INVCHD U536 ( .I(MK[32]), .O(n414) );
  NR2BHD U537 ( .I1(n148), .I2(n144), .O(n115) );
  INVCHD U538 ( .I(MK[0]), .O(n413) );
  OAI12CHD U539 ( .B1(n148), .B2(n149), .A1(n173), .O(n113) );
  ND2CHD U540 ( .I1(n162), .I2(n142), .O(n173) );
  NR3BHD U541 ( .I1(n579), .I2(n580), .I3(n581), .O(n162) );
  INVCHD U542 ( .I(MK[104]), .O(n303) );
  NR2BHD U543 ( .I1(n148), .I2(n93), .O(n153) );
  AO2222BHD U544 ( .A1(MK[112]), .A2(n27), .B1(MK[8]), .B2(n39), .C1(MK[40]), 
        .C2(n56), .D1(MK[72]), .D2(n143), .O(n575) );
  OAI12CHD U545 ( .B1(n578), .B2(n148), .A1(n174), .O(n143) );
  INVCHD U546 ( .I(n164), .O(n174) );
  NR2BHD U547 ( .I1(n109), .I2(n144), .O(n164) );
  INVCHD U548 ( .I(n123), .O(n148) );
  NR3BHD U549 ( .I1(n579), .I2(i_round[0]), .I3(n581), .O(n123) );
  OAI22CHD U550 ( .A1(n144), .A2(n145), .B1(n578), .B2(n109), .O(n189) );
  OAI22CHD U551 ( .A1(n149), .A2(n145), .B1(n93), .B2(n109), .O(n178) );
  INVCHD U552 ( .I(n582), .O(n109) );
  NR3BHD U553 ( .I1(n580), .I2(i_round[2]), .I3(n581), .O(n582) );
  INVCHD U554 ( .I(i_round[3]), .O(n581) );
  ND2CHD U555 ( .I1(n186), .I2(n141), .O(n106) );
  OA2222CHD U556 ( .A1(n126), .A2(n311), .B1(n118), .B2(n412), .C1(n32), .C2(
        n411), .D1(n120), .D2(n305), .O(n573) );
  INVCHD U557 ( .I(MK[80]), .O(n305) );
  ND2CHD U558 ( .I1(n133), .I2(n141), .O(n138) );
  ND3CHD U559 ( .I1(n580), .I2(n579), .I3(i_round[3]), .O(n145) );
  INVCHD U560 ( .I(MK[48]), .O(n411) );
  AN2CHD U561 ( .I1(n124), .I2(n141), .O(n152) );
  INVCHD U562 ( .I(MK[16]), .O(n412) );
  NR2BHD U563 ( .I1(n149), .I2(n156), .O(n159) );
  NR3BHD U564 ( .I1(n580), .I2(i_round[3]), .I3(n579), .O(n141) );
  INVCHD U565 ( .I(MK[120]), .O(n311) );
  NR2BHD U566 ( .I1(n171), .I2(n149), .O(n170) );
  AO2222BHD U567 ( .A1(mkx3[0]), .A2(n64), .B1(MK[24]), .B2(n188), .C1(MK[56]), 
        .C2(n38), .D1(MK[88]), .D2(n70), .O(n572) );
  INVCHD U568 ( .I(n136), .O(n206) );
  NR2BHD U569 ( .I1(n116), .I2(n166), .O(n136) );
  NR2BHD U570 ( .I1(n171), .I2(n144), .O(n166) );
  INVCHD U571 ( .I(n133), .O(n144) );
  NR2BHD U572 ( .I1(n156), .I2(n578), .O(n116) );
  INVCHD U573 ( .I(n124), .O(n578) );
  INVCHD U574 ( .I(n131), .O(n156) );
  NR3BHD U575 ( .I1(i_round[0]), .I2(i_round[3]), .I3(n579), .O(n131) );
  INVCHD U576 ( .I(i_round[2]), .O(n579) );
  INVCHD U577 ( .I(n134), .O(n177) );
  AOI22BHD U578 ( .A1(n132), .A2(n133), .B1(n124), .B2(n167), .O(n134) );
  NR3BHD U579 ( .I1(i_round[4]), .I2(i_round[5]), .I3(n584), .O(n133) );
  OAI12CHD U580 ( .B1(n93), .B2(n171), .A1(n150), .O(n188) );
  INVCHD U581 ( .I(n104), .O(n150) );
  NR2BHD U582 ( .I1(n149), .I2(n92), .O(n104) );
  INVCHD U583 ( .I(n186), .O(n149) );
  NR2BHD U584 ( .I1(n583), .I2(n584), .O(n186) );
  INVCHD U585 ( .I(i_round[1]), .O(n584) );
  INVCHD U586 ( .I(n167), .O(n171) );
  NR3BHD U587 ( .I1(i_round[2]), .I2(i_round[3]), .I3(n580), .O(n167) );
  INVCHD U588 ( .I(i_round[0]), .O(n580) );
  INVCHD U589 ( .I(n142), .O(n93) );
  NR2BHD U590 ( .I1(n91), .I2(i_round[5]), .O(n142) );
  INVCHD U591 ( .I(n585), .O(n91) );
  OA112CHD U592 ( .C1(n586), .C2(i_round[5]), .A1(n583), .B1(n187), .O(n205)
         );
  ND3CHD U593 ( .I1(n132), .I2(n585), .I3(i_round[5]), .O(n187) );
  NR2BHD U594 ( .I1(i_round[1]), .I2(i_round[4]), .O(n585) );
  OR2B1CHD U595 ( .I1(i_round[5]), .B1(i_round[4]), .O(n583) );
  NR2BHD U596 ( .I1(i_round[1]), .I2(n92), .O(n586) );
  INVCHD U597 ( .I(n132), .O(n92) );
  NR3BHD U598 ( .I1(i_round[2]), .I2(i_round[3]), .I3(i_round[0]), .O(n132) );
endmodule


module WK ( MK, clk, reset, ed, WK0_4, WK1_5, WK2_6, WK3_7 );
  input [127:0] MK;
  output [7:0] WK0_4;
  output [7:0] WK1_5;
  output [7:0] WK2_6;
  output [7:0] WK3_7;
  input clk, reset, ed;
  wire   MK_31, MK_30, MK_29, MK_28, MK_27, MK_26, MK_25, MK_24, MK_23, MK_22,
         MK_21, MK_20, MK_19, MK_18, MK_17, MK_16, MK_15, MK_14, MK_13, MK_12,
         MK_11, MK_10, MK_9, MK_8, MK_7, MK_6, MK_5, MK_4, MK_3, MK_2, MK_1,
         MK_0, N70, N71, N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N90, N91, N92, N93, N94, N95, N96,
         N97, N98, N99, N100, N101, N102, N105, N106, N107, N108, N109, n13,
         \add_32/carry[5] , \add_32/carry[4] , \add_32/carry[3] ,
         \add_32/carry[2] , n1, n2, n8, n9, n10;
  wire   [5:0] i_round;
  assign MK_31 = MK[31];
  assign MK_30 = MK[30];
  assign MK_29 = MK[29];
  assign MK_28 = MK[28];
  assign MK_27 = MK[27];
  assign MK_26 = MK[26];
  assign MK_25 = MK[25];
  assign MK_24 = MK[24];
  assign MK_23 = MK[23];
  assign MK_22 = MK[22];
  assign MK_21 = MK[21];
  assign MK_20 = MK[20];
  assign MK_19 = MK[19];
  assign MK_18 = MK[18];
  assign MK_17 = MK[17];
  assign MK_16 = MK[16];
  assign MK_15 = MK[15];
  assign MK_14 = MK[14];
  assign MK_13 = MK[13];
  assign MK_12 = MK[12];
  assign MK_11 = MK[11];
  assign MK_10 = MK[10];
  assign MK_9 = MK[9];
  assign MK_8 = MK[8];
  assign MK_7 = MK[7];
  assign MK_6 = MK[6];
  assign MK_5 = MK[5];
  assign MK_4 = MK[4];
  assign MK_3 = MK[3];
  assign MK_2 = MK[2];
  assign MK_1 = MK[1];
  assign MK_0 = MK[0];

  NR6EHD U39 ( .I1(i_round[3]), .I2(i_round[5]), .I3(i_round[4]), .I4(
        i_round[0]), .I5(i_round[2]), .I6(i_round[1]), .O(n13) );
  QDFFEHD \WK3_7_reg[5]  ( .D(N99), .CK(clk), .Q(WK3_7[5]) );
  QDFFEHD \WK3_7_reg[4]  ( .D(N98), .CK(clk), .Q(WK3_7[4]) );
  QDFFEHD \WK3_7_reg[3]  ( .D(N97), .CK(clk), .Q(WK3_7[3]) );
  QDFFEHD \WK3_7_reg[2]  ( .D(N96), .CK(clk), .Q(WK3_7[2]) );
  QDFFEHD \WK3_7_reg[1]  ( .D(N95), .CK(clk), .Q(WK3_7[1]) );
  QDFFEHD \WK3_7_reg[0]  ( .D(N94), .CK(clk), .Q(WK3_7[0]) );
  QDFFEHD \WK1_5_reg[7]  ( .D(N85), .CK(clk), .Q(WK1_5[7]) );
  QDFFEHD \WK1_5_reg[6]  ( .D(N84), .CK(clk), .Q(WK1_5[6]) );
  QDFFEHD \WK1_5_reg[5]  ( .D(N83), .CK(clk), .Q(WK1_5[5]) );
  QDFFEHD \WK1_5_reg[4]  ( .D(N82), .CK(clk), .Q(WK1_5[4]) );
  QDFFEHD \WK1_5_reg[3]  ( .D(N81), .CK(clk), .Q(WK1_5[3]) );
  QDFFEHD \WK1_5_reg[2]  ( .D(N80), .CK(clk), .Q(WK1_5[2]) );
  QDFFEHD \WK1_5_reg[1]  ( .D(N79), .CK(clk), .Q(WK1_5[1]) );
  QDFFEHD \WK1_5_reg[0]  ( .D(N78), .CK(clk), .Q(WK1_5[0]) );
  QDFFEHD \WK3_7_reg[7]  ( .D(N101), .CK(clk), .Q(WK3_7[7]) );
  QDFFEHD \WK3_7_reg[6]  ( .D(N100), .CK(clk), .Q(WK3_7[6]) );
  DFCLRBEHD \i_round_reg[5]  ( .RB(n10), .D(N109), .LD(N102), .CK(clk), .Q(
        i_round[5]) );
  DFCLRBEHD \i_round_reg[1]  ( .RB(n10), .D(N105), .LD(N102), .CK(clk), .Q(
        i_round[1]) );
  DFCLRBEHD \i_round_reg[2]  ( .RB(n10), .D(N106), .LD(N102), .CK(clk), .Q(
        i_round[2]) );
  DFCLRBEHD \i_round_reg[4]  ( .RB(n10), .D(N108), .LD(N102), .CK(clk), .Q(
        i_round[4]) );
  DFCLRBEHD \i_round_reg[3]  ( .RB(n10), .D(N107), .LD(N102), .CK(clk), .Q(
        i_round[3]) );
  DFCLRBEHD \i_round_reg[0]  ( .RB(n10), .D(n2), .LD(N102), .CK(clk), .Q(
        i_round[0]), .QB(n2) );
  QDFFEHD \WK2_6_reg[7]  ( .D(N93), .CK(clk), .Q(WK2_6[7]) );
  QDFFEHD \WK2_6_reg[6]  ( .D(N92), .CK(clk), .Q(WK2_6[6]) );
  QDFFEHD \WK2_6_reg[5]  ( .D(N91), .CK(clk), .Q(WK2_6[5]) );
  QDFFEHD \WK0_4_reg[7]  ( .D(N77), .CK(clk), .Q(WK0_4[7]) );
  QDFFEHD \WK0_4_reg[6]  ( .D(N76), .CK(clk), .Q(WK0_4[6]) );
  QDFFEHD \WK0_4_reg[5]  ( .D(N75), .CK(clk), .Q(WK0_4[5]) );
  QDFFEHD \WK2_6_reg[4]  ( .D(N90), .CK(clk), .Q(WK2_6[4]) );
  QDFFEHD \WK2_6_reg[3]  ( .D(N89), .CK(clk), .Q(WK2_6[3]) );
  QDFFEHD \WK2_6_reg[2]  ( .D(N88), .CK(clk), .Q(WK2_6[2]) );
  QDFFEHD \WK2_6_reg[1]  ( .D(N87), .CK(clk), .Q(WK2_6[1]) );
  QDFFEHD \WK2_6_reg[0]  ( .D(N86), .CK(clk), .Q(WK2_6[0]) );
  QDFFEHD \WK0_4_reg[4]  ( .D(N74), .CK(clk), .Q(WK0_4[4]) );
  QDFFEHD \WK0_4_reg[3]  ( .D(N73), .CK(clk), .Q(WK0_4[3]) );
  QDFFEHD \WK0_4_reg[2]  ( .D(N72), .CK(clk), .Q(WK0_4[2]) );
  QDFFEHD \WK0_4_reg[1]  ( .D(N71), .CK(clk), .Q(WK0_4[1]) );
  QDFFEHD \WK0_4_reg[0]  ( .D(N70), .CK(clk), .Q(WK0_4[0]) );
  XOR2EHD U3 ( .I1(ed), .I2(n13), .O(n1) );
  INVDHD U4 ( .I(n1), .O(n8) );
  AO22CHD U5 ( .A1(MK_30), .A2(n1), .B1(MK[126]), .B2(n8), .O(N100) );
  AO22CHD U6 ( .A1(MK_31), .A2(n1), .B1(MK[127]), .B2(n8), .O(N101) );
  AO22CHD U7 ( .A1(MK_0), .A2(n1), .B1(MK[96]), .B2(n8), .O(N70) );
  AO22CHD U8 ( .A1(MK_1), .A2(n1), .B1(MK[97]), .B2(n8), .O(N71) );
  AO22CHD U9 ( .A1(MK_2), .A2(n1), .B1(MK[98]), .B2(n8), .O(N72) );
  AO22CHD U10 ( .A1(MK_3), .A2(n1), .B1(MK[99]), .B2(n8), .O(N73) );
  AO22CHD U11 ( .A1(MK_4), .A2(n1), .B1(MK[100]), .B2(n8), .O(N74) );
  AO22CHD U12 ( .A1(MK_5), .A2(n1), .B1(MK[101]), .B2(n8), .O(N75) );
  AO22CHD U13 ( .A1(MK_6), .A2(n1), .B1(MK[102]), .B2(n8), .O(N76) );
  AO22CHD U14 ( .A1(MK_7), .A2(n1), .B1(MK[103]), .B2(n8), .O(N77) );
  AO22CHD U15 ( .A1(MK_8), .A2(n1), .B1(MK[104]), .B2(n8), .O(N78) );
  AO22CHD U16 ( .A1(MK_9), .A2(n1), .B1(MK[105]), .B2(n8), .O(N79) );
  AO22CHD U17 ( .A1(MK_10), .A2(n1), .B1(MK[106]), .B2(n8), .O(N80) );
  AO22CHD U18 ( .A1(MK_11), .A2(n1), .B1(MK[107]), .B2(n8), .O(N81) );
  AO22CHD U19 ( .A1(MK_12), .A2(n1), .B1(MK[108]), .B2(n8), .O(N82) );
  AO22CHD U20 ( .A1(MK_13), .A2(n1), .B1(MK[109]), .B2(n8), .O(N83) );
  AO22CHD U21 ( .A1(MK_14), .A2(n1), .B1(MK[110]), .B2(n8), .O(N84) );
  AO22CHD U22 ( .A1(MK_15), .A2(n1), .B1(MK[111]), .B2(n8), .O(N85) );
  AO22CHD U23 ( .A1(MK_16), .A2(n1), .B1(MK[112]), .B2(n8), .O(N86) );
  AO22CHD U24 ( .A1(MK_17), .A2(n1), .B1(MK[113]), .B2(n8), .O(N87) );
  AO22CHD U25 ( .A1(MK_18), .A2(n1), .B1(MK[114]), .B2(n8), .O(N88) );
  AO22CHD U26 ( .A1(MK_19), .A2(n1), .B1(MK[115]), .B2(n8), .O(N89) );
  AO22CHD U27 ( .A1(MK_20), .A2(n1), .B1(MK[116]), .B2(n8), .O(N90) );
  AO22CHD U28 ( .A1(MK_21), .A2(n1), .B1(MK[117]), .B2(n8), .O(N91) );
  AO22CHD U29 ( .A1(MK_22), .A2(n1), .B1(MK[118]), .B2(n8), .O(N92) );
  AO22CHD U30 ( .A1(MK_23), .A2(n1), .B1(MK[119]), .B2(n8), .O(N93) );
  AO22CHD U31 ( .A1(MK_24), .A2(n1), .B1(MK[120]), .B2(n8), .O(N94) );
  AO22CHD U32 ( .A1(MK_25), .A2(n1), .B1(MK[121]), .B2(n8), .O(N95) );
  AO22CHD U33 ( .A1(MK_26), .A2(n1), .B1(MK[122]), .B2(n8), .O(N96) );
  AO22CHD U34 ( .A1(MK_27), .A2(n1), .B1(MK[123]), .B2(n8), .O(N97) );
  AO22CHD U35 ( .A1(MK_28), .A2(n1), .B1(MK[124]), .B2(n8), .O(N98) );
  AO22CHD U36 ( .A1(MK_29), .A2(n1), .B1(MK[125]), .B2(n8), .O(N99) );
  INVDHD U37 ( .I(reset), .O(n10) );
  HA1EHD U38 ( .A(i_round[1]), .B(i_round[0]), .C(\add_32/carry[2] ), .S(N105)
         );
  HA1EHD U40 ( .A(i_round[3]), .B(\add_32/carry[3] ), .C(\add_32/carry[4] ), 
        .S(N107) );
  HA1EHD U41 ( .A(i_round[2]), .B(\add_32/carry[2] ), .C(\add_32/carry[3] ), 
        .S(N106) );
  HA1EHD U42 ( .A(i_round[4]), .B(\add_32/carry[4] ), .C(\add_32/carry[5] ), 
        .S(N108) );
  XOR2CHD U43 ( .I1(\add_32/carry[5] ), .I2(i_round[5]), .O(N109) );
  AO12CHD U44 ( .B1(i_round[1]), .B2(i_round[0]), .A1(i_round[2]), .O(n9) );
  OAI13BHD U45 ( .B1(n9), .B2(i_round[4]), .B3(i_round[3]), .A1(i_round[5]), 
        .O(N102) );
endmodule


module hight ( P, MK, clk, reset, ed, C );
  input [63:0] P;
  input [127:0] MK;
  output [63:0] C;
  input clk, reset, ed;

  wire   [7:0] WK0_4;
  wire   [7:0] WK1_5;
  wire   [7:0] WK2_6;
  wire   [7:0] WK3_7;
  wire   [7:0] SKx0;
  wire   [7:0] SKx1;
  wire   [7:0] SKx2;
  wire   [7:0] SKx3;

  WK whitening ( .MK(MK), .clk(clk), .reset(reset), .ed(ed), .WK0_4(WK0_4), 
        .WK1_5(WK1_5), .WK2_6(WK2_6), .WK3_7(WK3_7) );
  SK_gen subkey ( .MK(MK), .clk(clk), .reset(reset), .ed(ed), .SKx0(SKx0), 
        .SKx1(SKx1), .SKx2(SKx2), .SKx3(SKx3) );
  round_funct roundfunction ( .P(P), .MK(MK), .SKx0(SKx0), .SKx1(SKx1), .SKx2(
        SKx2), .SKx3(SKx3), .clk(clk), .reset(reset), .ed(ed), .WK0_4(WK0_4), 
        .WK1_5(WK1_5), .WK2_6(WK2_6), .WK3_7(WK3_7), .C(C) );
endmodule

