module NR6EHD (
	O, 
	I6, 
	I5, 
	I4, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I6;
   input I5;
   input I4;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module QDFFEHD (
	Q, 
	D, 
	CK, 
	GND, 
	VCC);
   output Q;
   input D;
   input CK;
   inout GND;
   inout VCC;
endmodule

module DFCLRBEHD (
	RB, 
	QB, 
	Q, 
	LD, 
	D, 
	CK, 
	GND, 
	VCC);
   input RB;
   output QB;
   output Q;
   input LD;
   input D;
   input CK;
   inout GND;
   inout VCC;
endmodule

module XOR2EHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module INVDHD (
	O, 
	I, 
	GND, 
	VCC);
   output O;
   input I;
   inout GND;
   inout VCC;
endmodule

module AO22CHD (
	O, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module HA1EHD (
	S, 
	C, 
	B, 
	A, 
	GND, 
	VCC);
   output S;
   output C;
   input B;
   input A;
   inout GND;
   inout VCC;
endmodule

module XOR2CHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module AO12CHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module OAI13BHD (
	O, 
	B3, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B3;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module FA1DHD (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	GND, 
	VCC);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout GND;
   inout VCC;
endmodule

module XOR3EHD (
	O, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module TIE0DHD (
	O, 
	GND, 
	VCC);
   output O;
   inout GND;
   inout VCC;
endmodule

module AOI12EHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AN2EHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module OA12EHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AO12EHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module NR2CHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module NR2BHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module AN2B1CHD (
	O, 
	I1, 
	B1, 
	GND, 
	VCC);
   output O;
   input I1;
   input B1;
   inout GND;
   inout VCC;
endmodule

module AO112CHD (
	O, 
	C2, 
	C1, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module MUX2CHD (
	S, 
	O, 
	B, 
	A, 
	GND, 
	VCC);
   input S;
   output O;
   input B;
   input A;
   inout GND;
   inout VCC;
endmodule

module OR3B2CHD (
	O, 
	I1, 
	B2, 
	B1, 
	GND, 
	VCC);
   output O;
   input I1;
   input B2;
   input B1;
   inout GND;
   inout VCC;
endmodule

module AOI22BHD (
	O, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AO222CHD (
	O, 
	C2, 
	C1, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module INVCHD (
	O, 
	I, 
	GND, 
	VCC);
   output O;
   input I;
   inout GND;
   inout VCC;
endmodule

module ND3CHD (
	O, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module ND2CHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module OAI12CHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module OAI112BHD (
	O, 
	C2, 
	C1, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AOI112BHD (
	O, 
	C2, 
	C1, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AN3B2BHD (
	O, 
	I1, 
	B2, 
	B1, 
	GND, 
	VCC);
   output O;
   input I1;
   input B2;
   input B1;
   inout GND;
   inout VCC;
endmodule

module ND6EHD (
	O, 
	I6, 
	I5, 
	I4, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I6;
   input I5;
   input I4;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module AN4B1BHD (
	O, 
	I3, 
	I2, 
	I1, 
	B1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   input B1;
   inout GND;
   inout VCC;
endmodule

module OA12CHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AOI12CHD (
	O, 
	B2, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module OA112CHD (
	O, 
	C2, 
	C1, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module NR3BHD (
	O, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module OAI22CHD (
	O, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module OAI222BHD (
	O, 
	C2, 
	C1, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AO2222BHD (
	O, 
	D2, 
	D1, 
	C2, 
	C1, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input D2;
   input D1;
   input C2;
   input C1;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module OA2222CHD (
	O, 
	D2, 
	D1, 
	C2, 
	C1, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input D2;
   input D1;
   input C2;
   input C1;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AN2CHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module OR2B1CHD (
	O, 
	I1, 
	B1, 
	GND, 
	VCC);
   output O;
   input I1;
   input B1;
   inout GND;
   inout VCC;
endmodule

module TIE1DHD (
	O, 
	GND, 
	VCC);
   output O;
   inout GND;
   inout VCC;
endmodule

module DFECHD (
	QB, 
	Q, 
	EB, 
	D, 
	CK, 
	GND, 
	VCC);
   output QB;
   output Q;
   input EB;
   input D;
   input CK;
   inout GND;
   inout VCC;
endmodule

module DFFCHD (
	QB, 
	Q, 
	D, 
	CK, 
	GND, 
	VCC);
   output QB;
   output Q;
   input D;
   input CK;
   inout GND;
   inout VCC;
endmodule

module AN3EHD (
	O, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module OA112EHD (
	O, 
	C2, 
	C1, 
	B1, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B1;
   input A1;
   inout GND;
   inout VCC;
endmodule

module AOI222BHD (
	O, 
	C2, 
	C1, 
	B2, 
	B1, 
	A2, 
	A1, 
	GND, 
	VCC);
   output O;
   input C2;
   input C1;
   input B2;
   input B1;
   input A2;
   input A1;
   inout GND;
   inout VCC;
endmodule

module ND2HHD (
	O, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module XOR4EHD (
	O, 
	I4, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I4;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module XOR3CHD (
	O, 
	I3, 
	I2, 
	I1, 
	GND, 
	VCC);
   output O;
   input I3;
   input I2;
   input I1;
   inout GND;
   inout VCC;
endmodule

module WK (
	MK, 
	clk, 
	reset, 
	ed, 
	WK0_4, 
	WK1_5, 
	WK2_6, 
	WK3_7);
   input [127:0] MK;
   input clk;
   input reset;
   input ed;
   output [7:0] WK0_4;
   output [7:0] WK1_5;
   output [7:0] WK2_6;
   output [7:0] WK3_7;

   // Internal wires
   wire MK_31;
   wire MK_30;
   wire MK_29;
   wire MK_28;
   wire MK_27;
   wire MK_26;
   wire MK_25;
   wire MK_24;
   wire MK_23;
   wire MK_22;
   wire MK_21;
   wire MK_20;
   wire MK_19;
   wire MK_18;
   wire MK_17;
   wire MK_16;
   wire MK_15;
   wire MK_14;
   wire MK_13;
   wire MK_12;
   wire MK_11;
   wire MK_10;
   wire MK_9;
   wire MK_8;
   wire MK_7;
   wire MK_6;
   wire MK_5;
   wire MK_4;
   wire MK_3;
   wire MK_2;
   wire MK_1;
   wire MK_0;
   wire N70;
   wire N71;
   wire N72;
   wire N73;
   wire N74;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire n13;
   wire \add_32/carry[5] ;
   wire \add_32/carry[4] ;
   wire \add_32/carry[3] ;
   wire \add_32/carry[2] ;
   wire n1;
   wire n2;
   wire n8;
   wire n9;
   wire n10;
   wire [5:0] i_round;

   assign MK_31 = MK[31] ;
   assign MK_30 = MK[30] ;
   assign MK_29 = MK[29] ;
   assign MK_28 = MK[28] ;
   assign MK_27 = MK[27] ;
   assign MK_26 = MK[26] ;
   assign MK_25 = MK[25] ;
   assign MK_24 = MK[24] ;
   assign MK_23 = MK[23] ;
   assign MK_22 = MK[22] ;
   assign MK_21 = MK[21] ;
   assign MK_20 = MK[20] ;
   assign MK_19 = MK[19] ;
   assign MK_18 = MK[18] ;
   assign MK_17 = MK[17] ;
   assign MK_16 = MK[16] ;
   assign MK_15 = MK[15] ;
   assign MK_14 = MK[14] ;
   assign MK_13 = MK[13] ;
   assign MK_12 = MK[12] ;
   assign MK_11 = MK[11] ;
   assign MK_10 = MK[10] ;
   assign MK_9 = MK[9] ;
   assign MK_8 = MK[8] ;
   assign MK_7 = MK[7] ;
   assign MK_6 = MK[6] ;
   assign MK_5 = MK[5] ;
   assign MK_4 = MK[4] ;
   assign MK_3 = MK[3] ;
   assign MK_2 = MK[2] ;
   assign MK_1 = MK[1] ;
   assign MK_0 = MK[0] ;

   // Module instantiations
   NR6EHD U39 (
	.O(n13),
	.I6(i_round[1]),
	.I5(i_round[2]),
	.I4(i_round[0]),
	.I3(i_round[4]),
	.I2(i_round[5]),
	.I1(i_round[3]));
   QDFFEHD \WK3_7_reg[5]  (
	.Q(WK3_7[5]),
	.D(N99),
	.CK(clk));
   QDFFEHD \WK3_7_reg[4]  (
	.Q(WK3_7[4]),
	.D(N98),
	.CK(clk));
   QDFFEHD \WK3_7_reg[3]  (
	.Q(WK3_7[3]),
	.D(N97),
	.CK(clk));
   QDFFEHD \WK3_7_reg[2]  (
	.Q(WK3_7[2]),
	.D(N96),
	.CK(clk));
   QDFFEHD \WK3_7_reg[1]  (
	.Q(WK3_7[1]),
	.D(N95),
	.CK(clk));
   QDFFEHD \WK3_7_reg[0]  (
	.Q(WK3_7[0]),
	.D(N94),
	.CK(clk));
   QDFFEHD \WK1_5_reg[7]  (
	.Q(WK1_5[7]),
	.D(N85),
	.CK(clk));
   QDFFEHD \WK1_5_reg[6]  (
	.Q(WK1_5[6]),
	.D(N84),
	.CK(clk));
   QDFFEHD \WK1_5_reg[5]  (
	.Q(WK1_5[5]),
	.D(N83),
	.CK(clk));
   QDFFEHD \WK1_5_reg[4]  (
	.Q(WK1_5[4]),
	.D(N82),
	.CK(clk));
   QDFFEHD \WK1_5_reg[3]  (
	.Q(WK1_5[3]),
	.D(N81),
	.CK(clk));
   QDFFEHD \WK1_5_reg[2]  (
	.Q(WK1_5[2]),
	.D(N80),
	.CK(clk));
   QDFFEHD \WK1_5_reg[1]  (
	.Q(WK1_5[1]),
	.D(N79),
	.CK(clk));
   QDFFEHD \WK1_5_reg[0]  (
	.Q(WK1_5[0]),
	.D(N78),
	.CK(clk));
   QDFFEHD \WK3_7_reg[7]  (
	.Q(WK3_7[7]),
	.D(N101),
	.CK(clk));
   QDFFEHD \WK3_7_reg[6]  (
	.Q(WK3_7[6]),
	.D(N100),
	.CK(clk));
   DFCLRBEHD \i_round_reg[5]  (
	.RB(n10),
	.Q(i_round[5]),
	.LD(N102),
	.D(N109),
	.CK(clk));
   DFCLRBEHD \i_round_reg[1]  (
	.RB(n10),
	.Q(i_round[1]),
	.LD(N102),
	.D(N105),
	.CK(clk));
   DFCLRBEHD \i_round_reg[2]  (
	.RB(n10),
	.Q(i_round[2]),
	.LD(N102),
	.D(N106),
	.CK(clk));
   DFCLRBEHD \i_round_reg[4]  (
	.RB(n10),
	.Q(i_round[4]),
	.LD(N102),
	.D(N108),
	.CK(clk));
   DFCLRBEHD \i_round_reg[3]  (
	.RB(n10),
	.Q(i_round[3]),
	.LD(N102),
	.D(N107),
	.CK(clk));
   DFCLRBEHD \i_round_reg[0]  (
	.RB(n10),
	.QB(n2),
	.Q(i_round[0]),
	.LD(N102),
	.D(n2),
	.CK(clk));
   QDFFEHD \WK2_6_reg[7]  (
	.Q(WK2_6[7]),
	.D(N93),
	.CK(clk));
   QDFFEHD \WK2_6_reg[6]  (
	.Q(WK2_6[6]),
	.D(N92),
	.CK(clk));
   QDFFEHD \WK2_6_reg[5]  (
	.Q(WK2_6[5]),
	.D(N91),
	.CK(clk));
   QDFFEHD \WK0_4_reg[7]  (
	.Q(WK0_4[7]),
	.D(N77),
	.CK(clk));
   QDFFEHD \WK0_4_reg[6]  (
	.Q(WK0_4[6]),
	.D(N76),
	.CK(clk));
   QDFFEHD \WK0_4_reg[5]  (
	.Q(WK0_4[5]),
	.D(N75),
	.CK(clk));
   QDFFEHD \WK2_6_reg[4]  (
	.Q(WK2_6[4]),
	.D(N90),
	.CK(clk));
   QDFFEHD \WK2_6_reg[3]  (
	.Q(WK2_6[3]),
	.D(N89),
	.CK(clk));
   QDFFEHD \WK2_6_reg[2]  (
	.Q(WK2_6[2]),
	.D(N88),
	.CK(clk));
   QDFFEHD \WK2_6_reg[1]  (
	.Q(WK2_6[1]),
	.D(N87),
	.CK(clk));
   QDFFEHD \WK2_6_reg[0]  (
	.Q(WK2_6[0]),
	.D(N86),
	.CK(clk));
   QDFFEHD \WK0_4_reg[4]  (
	.Q(WK0_4[4]),
	.D(N74),
	.CK(clk));
   QDFFEHD \WK0_4_reg[3]  (
	.Q(WK0_4[3]),
	.D(N73),
	.CK(clk));
   QDFFEHD \WK0_4_reg[2]  (
	.Q(WK0_4[2]),
	.D(N72),
	.CK(clk));
   QDFFEHD \WK0_4_reg[1]  (
	.Q(WK0_4[1]),
	.D(N71),
	.CK(clk));
   QDFFEHD \WK0_4_reg[0]  (
	.Q(WK0_4[0]),
	.D(N70),
	.CK(clk));
   XOR2EHD U3 (
	.O(n1),
	.I2(n13),
	.I1(ed));
   INVDHD U4 (
	.O(n8),
	.I(n1));
   AO22CHD U5 (
	.O(N100),
	.B2(n8),
	.B1(MK[126]),
	.A2(n1),
	.A1(MK_30));
   AO22CHD U6 (
	.O(N101),
	.B2(n8),
	.B1(MK[127]),
	.A2(n1),
	.A1(MK_31));
   AO22CHD U7 (
	.O(N70),
	.B2(n8),
	.B1(MK[96]),
	.A2(n1),
	.A1(MK_0));
   AO22CHD U8 (
	.O(N71),
	.B2(n8),
	.B1(MK[97]),
	.A2(n1),
	.A1(MK_1));
   AO22CHD U9 (
	.O(N72),
	.B2(n8),
	.B1(MK[98]),
	.A2(n1),
	.A1(MK_2));
   AO22CHD U10 (
	.O(N73),
	.B2(n8),
	.B1(MK[99]),
	.A2(n1),
	.A1(MK_3));
   AO22CHD U11 (
	.O(N74),
	.B2(n8),
	.B1(MK[100]),
	.A2(n1),
	.A1(MK_4));
   AO22CHD U12 (
	.O(N75),
	.B2(n8),
	.B1(MK[101]),
	.A2(n1),
	.A1(MK_5));
   AO22CHD U13 (
	.O(N76),
	.B2(n8),
	.B1(MK[102]),
	.A2(n1),
	.A1(MK_6));
   AO22CHD U14 (
	.O(N77),
	.B2(n8),
	.B1(MK[103]),
	.A2(n1),
	.A1(MK_7));
   AO22CHD U15 (
	.O(N78),
	.B2(n8),
	.B1(MK[104]),
	.A2(n1),
	.A1(MK_8));
   AO22CHD U16 (
	.O(N79),
	.B2(n8),
	.B1(MK[105]),
	.A2(n1),
	.A1(MK_9));
   AO22CHD U17 (
	.O(N80),
	.B2(n8),
	.B1(MK[106]),
	.A2(n1),
	.A1(MK_10));
   AO22CHD U18 (
	.O(N81),
	.B2(n8),
	.B1(MK[107]),
	.A2(n1),
	.A1(MK_11));
   AO22CHD U19 (
	.O(N82),
	.B2(n8),
	.B1(MK[108]),
	.A2(n1),
	.A1(MK_12));
   AO22CHD U20 (
	.O(N83),
	.B2(n8),
	.B1(MK[109]),
	.A2(n1),
	.A1(MK_13));
   AO22CHD U21 (
	.O(N84),
	.B2(n8),
	.B1(MK[110]),
	.A2(n1),
	.A1(MK_14));
   AO22CHD U22 (
	.O(N85),
	.B2(n8),
	.B1(MK[111]),
	.A2(n1),
	.A1(MK_15));
   AO22CHD U23 (
	.O(N86),
	.B2(n8),
	.B1(MK[112]),
	.A2(n1),
	.A1(MK_16));
   AO22CHD U24 (
	.O(N87),
	.B2(n8),
	.B1(MK[113]),
	.A2(n1),
	.A1(MK_17));
   AO22CHD U25 (
	.O(N88),
	.B2(n8),
	.B1(MK[114]),
	.A2(n1),
	.A1(MK_18));
   AO22CHD U26 (
	.O(N89),
	.B2(n8),
	.B1(MK[115]),
	.A2(n1),
	.A1(MK_19));
   AO22CHD U27 (
	.O(N90),
	.B2(n8),
	.B1(MK[116]),
	.A2(n1),
	.A1(MK_20));
   AO22CHD U28 (
	.O(N91),
	.B2(n8),
	.B1(MK[117]),
	.A2(n1),
	.A1(MK_21));
   AO22CHD U29 (
	.O(N92),
	.B2(n8),
	.B1(MK[118]),
	.A2(n1),
	.A1(MK_22));
   AO22CHD U30 (
	.O(N93),
	.B2(n8),
	.B1(MK[119]),
	.A2(n1),
	.A1(MK_23));
   AO22CHD U31 (
	.O(N94),
	.B2(n8),
	.B1(MK[120]),
	.A2(n1),
	.A1(MK_24));
   AO22CHD U32 (
	.O(N95),
	.B2(n8),
	.B1(MK[121]),
	.A2(n1),
	.A1(MK_25));
   AO22CHD U33 (
	.O(N96),
	.B2(n8),
	.B1(MK[122]),
	.A2(n1),
	.A1(MK_26));
   AO22CHD U34 (
	.O(N97),
	.B2(n8),
	.B1(MK[123]),
	.A2(n1),
	.A1(MK_27));
   AO22CHD U35 (
	.O(N98),
	.B2(n8),
	.B1(MK[124]),
	.A2(n1),
	.A1(MK_28));
   AO22CHD U36 (
	.O(N99),
	.B2(n8),
	.B1(MK[125]),
	.A2(n1),
	.A1(MK_29));
   INVDHD U37 (
	.O(n10),
	.I(reset));
   HA1EHD U38 (
	.S(N105),
	.C(\add_32/carry[2] ),
	.B(i_round[0]),
	.A(i_round[1]));
   HA1EHD U40 (
	.S(N107),
	.C(\add_32/carry[4] ),
	.B(\add_32/carry[3] ),
	.A(i_round[3]));
   HA1EHD U41 (
	.S(N106),
	.C(\add_32/carry[3] ),
	.B(\add_32/carry[2] ),
	.A(i_round[2]));
   HA1EHD U42 (
	.S(N108),
	.C(\add_32/carry[5] ),
	.B(\add_32/carry[4] ),
	.A(i_round[4]));
   XOR2CHD U43 (
	.O(N109),
	.I2(i_round[5]),
	.I1(\add_32/carry[5] ));
   AO12CHD U44 (
	.O(n9),
	.B2(i_round[0]),
	.B1(i_round[1]),
	.A1(i_round[2]));
   OAI13BHD U45 (
	.O(N102),
	.B3(i_round[3]),
	.B2(i_round[4]),
	.B1(n9),
	.A1(i_round[5]));
endmodule

module SK_gen_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module SK_gen_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module SK_gen_DW01_add_2 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module SK_gen_DW01_add_3 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module SK_gen (
	MK, 
	clk, 
	reset, 
	ed, 
	SKx0, 
	SKx1, 
	SKx2, 
	SKx3);
   input [127:0] MK;
   input clk;
   input reset;
   input ed;
   output [7:0] SKx0;
   output [7:0] SKx1;
   output [7:0] SKx2;
   output [7:0] SKx3;

   // Internal wires
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N89;
   wire N90;
   wire N91;
   wire N92;
   wire N93;
   wire n1;
   wire n478;
   wire n479;
   wire n480;
   wire n481;
   wire n482;
   wire n483;
   wire n484;
   wire n485;
   wire n486;
   wire n487;
   wire n488;
   wire n489;
   wire n490;
   wire n491;
   wire n492;
   wire n493;
   wire n494;
   wire n495;
   wire n496;
   wire n497;
   wire n498;
   wire n499;
   wire n500;
   wire n501;
   wire n502;
   wire n503;
   wire n504;
   wire n505;
   wire n506;
   wire n507;
   wire n508;
   wire n509;
   wire n510;
   wire n511;
   wire n512;
   wire n513;
   wire n514;
   wire n515;
   wire n516;
   wire n517;
   wire n518;
   wire n519;
   wire n520;
   wire n521;
   wire n522;
   wire n523;
   wire n524;
   wire n525;
   wire n526;
   wire n527;
   wire n528;
   wire n529;
   wire n530;
   wire n531;
   wire n532;
   wire n533;
   wire n534;
   wire n535;
   wire n536;
   wire n537;
   wire n538;
   wire n539;
   wire n540;
   wire n541;
   wire n542;
   wire n543;
   wire \add_35/carry[5] ;
   wire \add_35/carry[4] ;
   wire \add_35/carry[3] ;
   wire \add_35/carry[2] ;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n14;
   wire n27;
   wire n54;
   wire n55;
   wire n60;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n335;
   wire n336;
   wire n337;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n351;
   wire n352;
   wire n353;
   wire n354;
   wire n355;
   wire n356;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n367;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire n448;
   wire n449;
   wire n450;
   wire n451;
   wire n452;
   wire n453;
   wire n454;
   wire n455;
   wire n456;
   wire n457;
   wire n458;
   wire n459;
   wire n460;
   wire n461;
   wire n462;
   wire n463;
   wire n464;
   wire n465;
   wire n466;
   wire n467;
   wire n468;
   wire n469;
   wire n470;
   wire n471;
   wire n472;
   wire n473;
   wire n474;
   wire n475;
   wire n476;
   wire n477;
   wire n544;
   wire n545;
   wire n546;
   wire n547;
   wire n548;
   wire n549;
   wire n550;
   wire n551;
   wire n552;
   wire n553;
   wire n554;
   wire n555;
   wire n556;
   wire n557;
   wire n558;
   wire n559;
   wire n560;
   wire n561;
   wire n562;
   wire n563;
   wire n564;
   wire n565;
   wire n566;
   wire n567;
   wire n568;
   wire n569;
   wire n570;
   wire n571;
   wire n572;
   wire n573;
   wire n574;
   wire n575;
   wire n576;
   wire n577;
   wire n578;
   wire n579;
   wire n580;
   wire n581;
   wire n582;
   wire n583;
   wire n584;
   wire n585;
   wire n586;
   wire [5:0] i_round;
   wire [6:0] dx0;
   wire [6:0] dx1;
   wire [6:0] dx2;
   wire [6:0] dx3;
   wire [7:0] mkx0;
   wire [7:0] mkx1;
   wire [7:0] mkx2;
   wire [7:0] mkx3;

   // Module instantiations
   SK_gen_DW01_add_0 add_354 (
	.A({ mkx3[7],
		mkx3[6],
		mkx3[5],
		mkx3[4],
		mkx3[3],
		mkx3[2],
		mkx3[1],
		mkx3[0] }),
	.B({ n1,
		dx3[6],
		dx3[5],
		dx3[4],
		dx3[3],
		dx3[2],
		dx3[1],
		dx3[0] }),
	.CI(n1),
	.SUM({ SKx3[7],
		SKx3[6],
		SKx3[5],
		SKx3[4],
		SKx3[3],
		SKx3[2],
		SKx3[1],
		SKx3[0] }));
   SK_gen_DW01_add_1 add_353 (
	.A({ mkx2[7],
		mkx2[6],
		mkx2[5],
		mkx2[4],
		mkx2[3],
		mkx2[2],
		mkx2[1],
		mkx2[0] }),
	.B({ n1,
		dx2[6],
		dx2[5],
		dx2[4],
		dx2[3],
		dx2[2],
		dx2[1],
		dx2[0] }),
	.CI(n1),
	.SUM({ SKx2[7],
		SKx2[6],
		SKx2[5],
		SKx2[4],
		SKx2[3],
		SKx2[2],
		SKx2[1],
		SKx2[0] }));
   SK_gen_DW01_add_2 add_352 (
	.A({ mkx1[7],
		mkx1[6],
		mkx1[5],
		mkx1[4],
		mkx1[3],
		mkx1[2],
		mkx1[1],
		mkx1[0] }),
	.B({ n1,
		dx1[6],
		dx1[5],
		dx1[4],
		dx1[3],
		dx1[2],
		dx1[1],
		dx1[0] }),
	.CI(n1),
	.SUM({ SKx1[7],
		SKx1[6],
		SKx1[5],
		SKx1[4],
		SKx1[3],
		SKx1[2],
		SKx1[1],
		SKx1[0] }));
   SK_gen_DW01_add_3 add_351 (
	.A({ mkx0[7],
		mkx0[6],
		mkx0[5],
		mkx0[4],
		mkx0[3],
		mkx0[2],
		mkx0[1],
		mkx0[0] }),
	.B({ n1,
		dx0[6],
		dx0[5],
		dx0[4],
		dx0[3],
		dx0[2],
		dx0[1],
		dx0[0] }),
	.CI(n1),
	.SUM({ SKx0[7],
		SKx0[6],
		SKx0[5],
		SKx0[4],
		SKx0[3],
		SKx0[2],
		SKx0[1],
		SKx0[0] }));
   QDFFEHD \mkx0_reg[7]  (
	.Q(mkx0[7]),
	.D(n509),
	.CK(clk));
   QDFFEHD \mkx0_reg[6]  (
	.Q(mkx0[6]),
	.D(n508),
	.CK(clk));
   QDFFEHD \mkx0_reg[5]  (
	.Q(mkx0[5]),
	.D(n507),
	.CK(clk));
   QDFFEHD \mkx0_reg[4]  (
	.Q(mkx0[4]),
	.D(n506),
	.CK(clk));
   QDFFEHD \mkx0_reg[3]  (
	.Q(mkx0[3]),
	.D(n505),
	.CK(clk));
   QDFFEHD \mkx1_reg[7]  (
	.Q(mkx1[7]),
	.D(n501),
	.CK(clk));
   QDFFEHD \mkx1_reg[6]  (
	.Q(mkx1[6]),
	.D(n500),
	.CK(clk));
   QDFFEHD \mkx1_reg[5]  (
	.Q(mkx1[5]),
	.D(n499),
	.CK(clk));
   QDFFEHD \mkx1_reg[4]  (
	.Q(mkx1[4]),
	.D(n498),
	.CK(clk));
   QDFFEHD \mkx1_reg[3]  (
	.Q(mkx1[3]),
	.D(n497),
	.CK(clk));
   QDFFEHD \mkx1_reg[2]  (
	.Q(mkx1[2]),
	.D(n496),
	.CK(clk));
   QDFFEHD \mkx2_reg[7]  (
	.Q(mkx2[7]),
	.D(n493),
	.CK(clk));
   QDFFEHD \mkx2_reg[6]  (
	.Q(mkx2[6]),
	.D(n492),
	.CK(clk));
   QDFFEHD \mkx2_reg[5]  (
	.Q(mkx2[5]),
	.D(n491),
	.CK(clk));
   QDFFEHD \mkx2_reg[4]  (
	.Q(mkx2[4]),
	.D(n490),
	.CK(clk));
   QDFFEHD \mkx2_reg[3]  (
	.Q(mkx2[3]),
	.D(n489),
	.CK(clk));
   QDFFEHD \mkx3_reg[7]  (
	.Q(mkx3[7]),
	.D(n485),
	.CK(clk));
   QDFFEHD \mkx3_reg[6]  (
	.Q(mkx3[6]),
	.D(n484),
	.CK(clk));
   QDFFEHD \mkx3_reg[5]  (
	.Q(mkx3[5]),
	.D(n483),
	.CK(clk));
   QDFFEHD \mkx3_reg[4]  (
	.Q(mkx3[4]),
	.D(n482),
	.CK(clk));
   QDFFEHD \mkx3_reg[3]  (
	.Q(mkx3[3]),
	.D(n481),
	.CK(clk));
   QDFFEHD \mkx3_reg[2]  (
	.Q(mkx3[2]),
	.D(n480),
	.CK(clk));
   QDFFEHD \dx0_reg[6]  (
	.Q(dx0[6]),
	.D(n537),
	.CK(clk));
   QDFFEHD \dx0_reg[5]  (
	.Q(dx0[5]),
	.D(n536),
	.CK(clk));
   QDFFEHD \dx0_reg[4]  (
	.Q(dx0[4]),
	.D(n535),
	.CK(clk));
   QDFFEHD \dx0_reg[3]  (
	.Q(dx0[3]),
	.D(n534),
	.CK(clk));
   QDFFEHD \dx1_reg[6]  (
	.Q(dx1[6]),
	.D(n530),
	.CK(clk));
   QDFFEHD \dx1_reg[5]  (
	.Q(dx1[5]),
	.D(n529),
	.CK(clk));
   QDFFEHD \dx1_reg[4]  (
	.Q(dx1[4]),
	.D(n528),
	.CK(clk));
   QDFFEHD \dx1_reg[3]  (
	.Q(dx1[3]),
	.D(n527),
	.CK(clk));
   QDFFEHD \dx1_reg[2]  (
	.Q(dx1[2]),
	.D(n526),
	.CK(clk));
   QDFFEHD \dx2_reg[6]  (
	.Q(dx2[6]),
	.D(n523),
	.CK(clk));
   QDFFEHD \dx2_reg[5]  (
	.Q(dx2[5]),
	.D(n522),
	.CK(clk));
   QDFFEHD \dx2_reg[4]  (
	.Q(dx2[4]),
	.D(n521),
	.CK(clk));
   QDFFEHD \dx2_reg[3]  (
	.Q(dx2[3]),
	.D(n520),
	.CK(clk));
   QDFFEHD \dx3_reg[5]  (
	.Q(dx3[5]),
	.D(n515),
	.CK(clk));
   QDFFEHD \dx3_reg[4]  (
	.Q(dx3[4]),
	.D(n514),
	.CK(clk));
   QDFFEHD \dx3_reg[3]  (
	.Q(dx3[3]),
	.D(n513),
	.CK(clk));
   QDFFEHD \dx3_reg[2]  (
	.Q(dx3[2]),
	.D(n512),
	.CK(clk));
   QDFFEHD \dx3_reg[6]  (
	.Q(dx3[6]),
	.D(n516),
	.CK(clk));
   QDFFEHD \mkx0_reg[2]  (
	.Q(mkx0[2]),
	.D(n504),
	.CK(clk));
   QDFFEHD \mkx0_reg[1]  (
	.Q(mkx0[1]),
	.D(n503),
	.CK(clk));
   QDFFEHD \mkx0_reg[0]  (
	.Q(mkx0[0]),
	.D(n502),
	.CK(clk));
   QDFFEHD \mkx1_reg[1]  (
	.Q(mkx1[1]),
	.D(n495),
	.CK(clk));
   QDFFEHD \mkx1_reg[0]  (
	.Q(mkx1[0]),
	.D(n494),
	.CK(clk));
   QDFFEHD \mkx2_reg[2]  (
	.Q(mkx2[2]),
	.D(n488),
	.CK(clk));
   QDFFEHD \mkx2_reg[1]  (
	.Q(mkx2[1]),
	.D(n487),
	.CK(clk));
   QDFFEHD \mkx2_reg[0]  (
	.Q(mkx2[0]),
	.D(n486),
	.CK(clk));
   QDFFEHD \mkx3_reg[1]  (
	.Q(mkx3[1]),
	.D(n479),
	.CK(clk));
   QDFFEHD \mkx3_reg[0]  (
	.Q(mkx3[0]),
	.D(n478),
	.CK(clk));
   QDFFEHD \dx0_reg[2]  (
	.Q(dx0[2]),
	.D(n533),
	.CK(clk));
   QDFFEHD \dx0_reg[1]  (
	.Q(dx0[1]),
	.D(n532),
	.CK(clk));
   QDFFEHD \dx1_reg[1]  (
	.Q(dx1[1]),
	.D(n525),
	.CK(clk));
   QDFFEHD \dx1_reg[0]  (
	.Q(dx1[0]),
	.D(n524),
	.CK(clk));
   QDFFEHD \dx2_reg[2]  (
	.Q(dx2[2]),
	.D(n519),
	.CK(clk));
   QDFFEHD \dx2_reg[1]  (
	.Q(dx2[1]),
	.D(n518),
	.CK(clk));
   QDFFEHD \dx2_reg[0]  (
	.Q(dx2[0]),
	.D(n517),
	.CK(clk));
   QDFFEHD \dx3_reg[1]  (
	.Q(dx3[1]),
	.D(n511),
	.CK(clk));
   QDFFEHD \dx3_reg[0]  (
	.Q(dx3[0]),
	.D(n510),
	.CK(clk));
   QDFFEHD \dx0_reg[0]  (
	.Q(dx0[0]),
	.D(n531),
	.CK(clk));
   QDFFEHD \i_round_reg[3]  (
	.Q(i_round[3]),
	.D(n539),
	.CK(clk));
   QDFFEHD \i_round_reg[4]  (
	.Q(i_round[4]),
	.D(n538),
	.CK(clk));
   QDFFEHD \i_round_reg[5]  (
	.Q(i_round[5]),
	.D(n542),
	.CK(clk));
   QDFFEHD \i_round_reg[2]  (
	.Q(i_round[2]),
	.D(n540),
	.CK(clk));
   QDFFEHD \i_round_reg[0]  (
	.Q(i_round[0]),
	.D(n543),
	.CK(clk));
   QDFFEHD \i_round_reg[1]  (
	.Q(i_round[1]),
	.D(n541),
	.CK(clk));
   AOI12EHD U3 (
	.O(n2),
	.B2(n162),
	.B1(n124),
	.A1(n115));
   AOI12EHD U4 (
	.O(n3),
	.B2(n186),
	.B1(n582),
	.A1(n153));
   AOI12EHD U5 (
	.O(n4),
	.B2(n133),
	.B1(n131),
	.A1(n152));
   AOI12EHD U6 (
	.O(n5),
	.B2(n186),
	.B1(n162),
	.A1(n140));
   AOI12EHD U7 (
	.O(n6),
	.B2(n162),
	.B1(n133),
	.A1(n158));
   INVDHD U19 (
	.O(n27),
	.I(n7));
   INVDHD U23 (
	.O(n54),
	.I(n188));
   INVDHD U25 (
	.O(n121),
	.I(n113));
   INVDHD U27 (
	.O(n14),
	.I(n143));
   INVDHD U28 (
	.O(n55),
	.I(n60));
   INVDHD U50 (
	.O(n60),
	.I(n189));
   AOI12EHD U70 (
	.O(n118),
	.B2(n141),
	.B1(n142),
	.A1(n159));
   AN2EHD U71 (
	.O(n94),
	.I2(n180),
	.I1(n179));
   OA12EHD U72 (
	.O(n7),
	.B2(n145),
	.B1(n93),
	.A1(n106));
   AO12EHD U73 (
	.O(n8),
	.B2(n131),
	.B1(n142),
	.A1(n170));
   INVDHD U74 (
	.O(n126),
	.I(n8));
   INVDHD U76 (
	.O(n77),
	.I(n73));
   INVDHD U77 (
	.O(n78),
	.I(n74));
   NR2CHD U80 (
	.O(n124),
	.I2(i_round[1]),
	.I1(n583));
   HA1EHD U81 (
	.S(N75),
	.C(\add_35/carry[2] ),
	.B(i_round[0]),
	.A(i_round[1]));
   HA1EHD U82 (
	.S(N76),
	.C(\add_35/carry[3] ),
	.B(\add_35/carry[2] ),
	.A(i_round[2]));
   HA1EHD U83 (
	.S(N77),
	.C(\add_35/carry[4] ),
	.B(\add_35/carry[3] ),
	.A(i_round[3]));
   HA1EHD U84 (
	.S(N78),
	.C(\add_35/carry[5] ),
	.B(\add_35/carry[4] ),
	.A(i_round[4]));
   TIE0DHD U85 (
	.O(n1));
   OA12EHD U86 (
	.O(n120),
	.B2(n145),
	.B1(n578),
	.A1(n138));
   XOR2CHD U87 (
	.O(N79),
	.I2(i_round[5]),
	.I1(\add_35/carry[5] ));
   NR2BHD U88 (
	.O(n73),
	.I2(i_round[0]),
	.I1(i_round[1]));
   AO12CHD U89 (
	.O(N89),
	.B2(i_round[1]),
	.B1(i_round[0]),
	.A1(n73));
   NR2BHD U90 (
	.O(n74),
	.I2(i_round[2]),
	.I1(n77));
   AO12CHD U91 (
	.O(N90),
	.B2(i_round[2]),
	.B1(n77),
	.A1(n74));
   NR2BHD U92 (
	.O(n75),
	.I2(i_round[3]),
	.I1(n78));
   AO12CHD U93 (
	.O(N91),
	.B2(i_round[3]),
	.B1(n78),
	.A1(n75));
   XOR2CHD U94 (
	.O(N92),
	.I2(n75),
	.I1(i_round[4]));
   AN2B1CHD U95 (
	.O(n76),
	.I1(n75),
	.B1(i_round[4]));
   XOR2CHD U96 (
	.O(N93),
	.I2(n76),
	.I1(i_round[5]));
   AO112CHD U97 (
	.O(n543),
	.C2(n79),
	.C1(n580),
	.B1(n81),
	.A1(n80));
   MUX2CHD U98 (
	.S(i_round[0]),
	.O(n81),
	.B(n83),
	.A(n82));
   OR3B2CHD U99 (
	.O(n542),
	.I1(n80),
	.B2(n85),
	.B1(n84));
   AOI22BHD U100 (
	.O(n85),
	.B2(n82),
	.B1(N79),
	.A2(n79),
	.A1(N93));
   NR2BHD U101 (
	.O(n80),
	.I2(ed),
	.I1(n86));
   AO222CHD U102 (
	.O(n541),
	.C2(n82),
	.C1(N75),
	.B2(n83),
	.B1(i_round[1]),
	.A2(n79),
	.A1(N89));
   AO222CHD U103 (
	.O(n540),
	.C2(n82),
	.C1(N76),
	.B2(n83),
	.B1(i_round[2]),
	.A2(n79),
	.A1(N90));
   AO222CHD U104 (
	.O(n539),
	.C2(n82),
	.C1(N77),
	.B2(n83),
	.B1(i_round[3]),
	.A2(n79),
	.A1(N91));
   AO222CHD U105 (
	.O(n538),
	.C2(n82),
	.C1(N78),
	.B2(n83),
	.B1(i_round[4]),
	.A2(n79),
	.A1(N92));
   NR2BHD U106 (
	.O(n82),
	.I2(n88),
	.I1(n87));
   INVCHD U107 (
	.O(n83),
	.I(n84));
   ND3CHD U108 (
	.O(n84),
	.I3(n89),
	.I2(n86),
	.I1(n88));
   ND2CHD U109 (
	.O(n88),
	.I2(n86),
	.I1(n90));
   OAI12CHD U110 (
	.O(n90),
	.B2(n92),
	.B1(n91),
	.A1(i_round[5]));
   INVCHD U111 (
	.O(n79),
	.I(n89));
   OAI112BHD U112 (
	.O(n89),
	.C2(n92),
	.C1(n93),
	.B1(n86),
	.A1(n87));
   INVCHD U113 (
	.O(n86),
	.I(reset));
   INVCHD U114 (
	.O(n87),
	.I(ed));
   AO12CHD U115 (
	.O(n537),
	.B2(n94),
	.B1(dx0[6]),
	.A1(n95));
   AO12CHD U116 (
	.O(n536),
	.B2(n94),
	.B1(dx0[5]),
	.A1(n96));
   AO12CHD U117 (
	.O(n535),
	.B2(n94),
	.B1(dx0[4]),
	.A1(n97));
   AO12CHD U118 (
	.O(n534),
	.B2(n94),
	.B1(dx0[3]),
	.A1(n98));
   AO12CHD U119 (
	.O(n533),
	.B2(n94),
	.B1(dx0[2]),
	.A1(n99));
   AO12CHD U120 (
	.O(n532),
	.B2(n94),
	.B1(dx0[1]),
	.A1(n100));
   OR3B2CHD U121 (
	.O(n531),
	.I1(n101),
	.B2(n103),
	.B1(n102));
   AOI112BHD U122 (
	.O(n103),
	.C2(n94),
	.C1(dx0[0]),
	.B1(n105),
	.A1(n104));
   INVCHD U123 (
	.O(n105),
	.I(n106));
   AO12CHD U124 (
	.O(n530),
	.B2(n94),
	.B1(dx1[6]),
	.A1(n107));
   AO12CHD U125 (
	.O(n529),
	.B2(n94),
	.B1(dx1[5]),
	.A1(n95));
   AO12CHD U126 (
	.O(n528),
	.B2(n94),
	.B1(dx1[4]),
	.A1(n96));
   AO12CHD U127 (
	.O(n527),
	.B2(n94),
	.B1(dx1[3]),
	.A1(n97));
   AO12CHD U128 (
	.O(n526),
	.B2(n94),
	.B1(dx1[2]),
	.A1(n98));
   AO12CHD U129 (
	.O(n525),
	.B2(n94),
	.B1(dx1[1]),
	.A1(n99));
   AO12CHD U130 (
	.O(n524),
	.B2(n94),
	.B1(dx1[0]),
	.A1(n100));
   OAI112BHD U131 (
	.O(n100),
	.C2(n109),
	.C1(n108),
	.B1(n111),
	.A1(n110));
   AN3B2BHD U132 (
	.O(n111),
	.I1(n112),
	.B2(n114),
	.B1(n113));
   NR2BHD U133 (
	.O(n110),
	.I2(n116),
	.I1(n115));
   AO12CHD U134 (
	.O(n523),
	.B2(n94),
	.B1(dx2[6]),
	.A1(n117));
   AO12CHD U135 (
	.O(n522),
	.B2(n94),
	.B1(dx2[5]),
	.A1(n107));
   AO12CHD U136 (
	.O(n521),
	.B2(n94),
	.B1(dx2[4]),
	.A1(n95));
   AO12CHD U137 (
	.O(n520),
	.B2(n94),
	.B1(dx2[3]),
	.A1(n96));
   AO12CHD U138 (
	.O(n519),
	.B2(n94),
	.B1(dx2[2]),
	.A1(n97));
   AO12CHD U139 (
	.O(n518),
	.B2(n94),
	.B1(dx2[1]),
	.A1(n98));
   AO12CHD U140 (
	.O(n517),
	.B2(n94),
	.B1(dx2[0]),
	.A1(n99));
   ND6EHD U141 (
	.O(n99),
	.I6(n122),
	.I5(n121),
	.I4(n120),
	.I3(n119),
	.I2(n118),
	.I1(n7));
   AOI112BHD U142 (
	.O(n122),
	.C2(n124),
	.C1(n123),
	.B1(n8),
	.A1(n125));
   OAI112BHD U143 (
	.O(n125),
	.C2(n128),
	.C1(n127),
	.B1(n130),
	.A1(n129));
   INVCHD U144 (
	.O(n130),
	.I(n116));
   OAI12CHD U145 (
	.O(n129),
	.B2(n132),
	.B1(n131),
	.A1(n133));
   ND6EHD U146 (
	.O(n516),
	.I6(n137),
	.I5(n14),
	.I4(n136),
	.I3(n135),
	.I2(n134),
	.I1(n119));
   AN4B1BHD U147 (
	.O(n137),
	.I3(n139),
	.I2(n138),
	.I1(n106),
	.B1(n140));
   AOI22BHD U148 (
	.O(n139),
	.B2(n142),
	.B1(n141),
	.A2(n94),
	.A1(dx3[6]));
   OA12CHD U149 (
	.O(n119),
	.B2(n145),
	.B1(n144),
	.A1(n6));
   AO12CHD U150 (
	.O(n515),
	.B2(n94),
	.B1(dx3[5]),
	.A1(n117));
   ND6EHD U151 (
	.O(n117),
	.I6(n147),
	.I5(n146),
	.I4(n5),
	.I3(n135),
	.I2(n7),
	.I1(n120));
   AOI12CHD U152 (
	.O(n147),
	.B2(n142),
	.B1(n131),
	.A1(n115));
   OA112CHD U153 (
	.O(n135),
	.C2(n149),
	.C1(n148),
	.B1(n151),
	.A1(n150));
   NR2BHD U154 (
	.O(n151),
	.I2(n153),
	.I1(n152));
   AO12CHD U155 (
	.O(n514),
	.B2(n94),
	.B1(dx3[4]),
	.A1(n107));
   OAI112BHD U156 (
	.O(n107),
	.C2(n145),
	.C1(n93),
	.B1(n154),
	.A1(n54));
   NR2BHD U157 (
	.O(n154),
	.I2(n101),
	.I1(n155));
   OAI112BHD U158 (
	.O(n101),
	.C2(n144),
	.C1(n156),
	.B1(n157),
	.A1(n60));
   NR3BHD U159 (
	.O(n157),
	.I3(n159),
	.I2(n158),
	.I1(n140));
   AO12CHD U160 (
	.O(n513),
	.B2(n94),
	.B1(dx3[3]),
	.A1(n95));
   AO12CHD U161 (
	.O(n512),
	.B2(n94),
	.B1(dx3[2]),
	.A1(n96));
   ND6EHD U162 (
	.O(n96),
	.I6(n161),
	.I5(n112),
	.I4(n5),
	.I3(n160),
	.I2(n126),
	.I1(n4));
   AOI112BHD U163 (
	.O(n161),
	.C2(n124),
	.C1(n162),
	.B1(n164),
	.A1(n163));
   OR3B2CHD U164 (
	.O(n163),
	.I1(n159),
	.B2(n150),
	.B1(n165));
   INVCHD U165 (
	.O(n165),
	.I(n166));
   AOI12CHD U166 (
	.O(n112),
	.B2(n167),
	.B1(n124),
	.A1(n153));
   AO12CHD U167 (
	.O(n511),
	.B2(n94),
	.B1(dx3[1]),
	.A1(n97));
   ND6EHD U168 (
	.O(n97),
	.I6(n169),
	.I5(n168),
	.I4(n118),
	.I3(n6),
	.I2(n160),
	.I1(n5));
   NR2BHD U169 (
	.O(n169),
	.I2(n152),
	.I1(n170));
   AO12CHD U170 (
	.O(n168),
	.B2(n171),
	.B1(n109),
	.A1(n108));
   AO12CHD U171 (
	.O(n510),
	.B2(n94),
	.B1(dx3[0]),
	.A1(n98));
   OAI112BHD U172 (
	.O(n98),
	.C2(n171),
	.C1(n93),
	.B1(n172),
	.A1(n102));
   NR2BHD U173 (
	.O(n172),
	.I2(n27),
	.I1(n155));
   ND3CHD U174 (
	.O(n155),
	.I3(n175),
	.I2(n174),
	.I1(n173));
   AN3B2BHD U175 (
	.O(n175),
	.I1(n138),
	.B2(n153),
	.B1(n170));
   AN3B2BHD U176 (
	.O(n102),
	.I1(n176),
	.B2(n115),
	.B1(n116));
   NR2BHD U177 (
	.O(n176),
	.I2(n178),
	.I1(n177));
   NR3BHD U178 (
	.O(n180),
	.I3(n140),
	.I2(n164),
	.I1(n181));
   OAI12CHD U179 (
	.O(n181),
	.B2(n145),
	.B1(n149),
	.A1(n160));
   OA12CHD U180 (
	.O(n160),
	.B2(n145),
	.B1(n108),
	.A1(n173));
   NR2BHD U181 (
	.O(n108),
	.I2(n124),
	.I1(n142));
   AN4B1BHD U182 (
	.O(n179),
	.I3(n134),
	.I2(n146),
	.I1(n60),
	.B1(n95));
   ND2CHD U183 (
	.O(n95),
	.I2(n183),
	.I1(n182));
   AOI112BHD U184 (
	.O(n183),
	.C2(n184),
	.C1(n123),
	.B1(n166),
	.A1(n185));
   OAI22CHD U185 (
	.O(n185),
	.B2(n149),
	.B1(n128),
	.A2(n109),
	.A1(n93));
   INVCHD U186 (
	.O(n128),
	.I(n162));
   INVCHD U187 (
	.O(n184),
	.I(n127));
   NR2BHD U188 (
	.O(n127),
	.I2(n124),
	.I1(n186));
   AN4B1BHD U189 (
	.O(n182),
	.I3(n3),
	.I2(n2),
	.I1(n4),
	.B1(n114));
   ND6EHD U190 (
	.O(n114),
	.I6(n106),
	.I5(n187),
	.I4(n138),
	.I3(n54),
	.I2(n126),
	.I1(n118));
   AOI12CHD U191 (
	.O(n146),
	.B2(n162),
	.B1(n133),
	.A1(n116));
   OR3B2CHD U192 (
	.O(n509),
	.I1(n190),
	.B2(n192),
	.B1(n191));
   NR3BHD U193 (
	.O(n192),
	.I3(n195),
	.I2(n194),
	.I1(n193));
   OAI22CHD U194 (
	.O(n195),
	.B2(n197),
	.B1(n5),
	.A2(n196),
	.A1(n6));
   OAI222BHD U195 (
	.O(n194),
	.C2(n200),
	.C1(n2),
	.B2(n199),
	.B1(n121),
	.A2(n198),
	.A1(n3));
   AO2222BHD U196 (
	.O(n193),
	.D2(n143),
	.D1(MK[119]),
	.C2(n55),
	.C1(MK[23]),
	.B2(n178),
	.B1(MK[55]),
	.A2(n27),
	.A1(MK[95]));
   OA2222CHD U197 (
	.O(n191),
	.D2(n204),
	.D1(n120),
	.C2(n203),
	.C1(n4),
	.B2(n202),
	.B1(n118),
	.A2(n201),
	.A1(n126));
   AO2222BHD U198 (
	.O(n190),
	.D2(n206),
	.D1(MK[71]),
	.C2(n177),
	.C1(MK[39]),
	.B2(n188),
	.B1(MK[7]),
	.A2(n205),
	.A1(mkx0[7]));
   OR3B2CHD U199 (
	.O(n508),
	.I1(n207),
	.B2(n209),
	.B1(n208));
   NR3BHD U200 (
	.O(n209),
	.I3(n212),
	.I2(n211),
	.I1(n210));
   OAI22CHD U201 (
	.O(n212),
	.B2(n214),
	.B1(n5),
	.A2(n213),
	.A1(n6));
   OAI222BHD U202 (
	.O(n211),
	.C2(n217),
	.C1(n2),
	.B2(n216),
	.B1(n121),
	.A2(n215),
	.A1(n3));
   AO2222BHD U203 (
	.O(n210),
	.D2(n143),
	.D1(MK[118]),
	.C2(n55),
	.C1(MK[22]),
	.B2(n178),
	.B1(MK[54]),
	.A2(n27),
	.A1(MK[94]));
   OA2222CHD U204 (
	.O(n208),
	.D2(n221),
	.D1(n120),
	.C2(n220),
	.C1(n4),
	.B2(n219),
	.B1(n118),
	.A2(n218),
	.A1(n126));
   AO2222BHD U205 (
	.O(n207),
	.D2(n206),
	.D1(MK[70]),
	.C2(n177),
	.C1(MK[38]),
	.B2(n188),
	.B1(MK[6]),
	.A2(n205),
	.A1(mkx0[6]));
   OR3B2CHD U206 (
	.O(n507),
	.I1(n222),
	.B2(n224),
	.B1(n223));
   NR3BHD U207 (
	.O(n224),
	.I3(n227),
	.I2(n226),
	.I1(n225));
   OAI22CHD U208 (
	.O(n227),
	.B2(n229),
	.B1(n5),
	.A2(n228),
	.A1(n6));
   OAI222BHD U209 (
	.O(n226),
	.C2(n232),
	.C1(n2),
	.B2(n231),
	.B1(n121),
	.A2(n230),
	.A1(n3));
   AO2222BHD U210 (
	.O(n225),
	.D2(n143),
	.D1(MK[117]),
	.C2(n55),
	.C1(MK[21]),
	.B2(n178),
	.B1(MK[53]),
	.A2(n27),
	.A1(MK[93]));
   OA2222CHD U211 (
	.O(n223),
	.D2(n236),
	.D1(n120),
	.C2(n235),
	.C1(n4),
	.B2(n234),
	.B1(n118),
	.A2(n233),
	.A1(n126));
   AO2222BHD U212 (
	.O(n222),
	.D2(n206),
	.D1(MK[69]),
	.C2(n177),
	.C1(MK[37]),
	.B2(n188),
	.B1(MK[5]),
	.A2(n205),
	.A1(mkx0[5]));
   OR3B2CHD U213 (
	.O(n506),
	.I1(n237),
	.B2(n239),
	.B1(n238));
   NR3BHD U214 (
	.O(n239),
	.I3(n242),
	.I2(n241),
	.I1(n240));
   OAI22CHD U215 (
	.O(n242),
	.B2(n244),
	.B1(n5),
	.A2(n243),
	.A1(n6));
   OAI222BHD U216 (
	.O(n241),
	.C2(n247),
	.C1(n2),
	.B2(n246),
	.B1(n121),
	.A2(n245),
	.A1(n3));
   AO2222BHD U217 (
	.O(n240),
	.D2(n143),
	.D1(MK[116]),
	.C2(n55),
	.C1(MK[20]),
	.B2(n178),
	.B1(MK[52]),
	.A2(n27),
	.A1(MK[92]));
   OA2222CHD U218 (
	.O(n238),
	.D2(n251),
	.D1(n120),
	.C2(n250),
	.C1(n4),
	.B2(n249),
	.B1(n118),
	.A2(n248),
	.A1(n126));
   AO2222BHD U219 (
	.O(n237),
	.D2(n206),
	.D1(MK[68]),
	.C2(n177),
	.C1(MK[36]),
	.B2(n188),
	.B1(MK[4]),
	.A2(n205),
	.A1(mkx0[4]));
   OR3B2CHD U220 (
	.O(n505),
	.I1(n252),
	.B2(n254),
	.B1(n253));
   NR3BHD U221 (
	.O(n254),
	.I3(n257),
	.I2(n256),
	.I1(n255));
   OAI22CHD U222 (
	.O(n257),
	.B2(n259),
	.B1(n5),
	.A2(n258),
	.A1(n6));
   OAI222BHD U223 (
	.O(n256),
	.C2(n262),
	.C1(n2),
	.B2(n261),
	.B1(n121),
	.A2(n260),
	.A1(n3));
   AO2222BHD U224 (
	.O(n255),
	.D2(n143),
	.D1(MK[115]),
	.C2(n55),
	.C1(MK[19]),
	.B2(n178),
	.B1(MK[51]),
	.A2(n27),
	.A1(MK[91]));
   OA2222CHD U225 (
	.O(n253),
	.D2(n266),
	.D1(n120),
	.C2(n265),
	.C1(n4),
	.B2(n264),
	.B1(n118),
	.A2(n263),
	.A1(n126));
   AO2222BHD U226 (
	.O(n252),
	.D2(n206),
	.D1(MK[67]),
	.C2(n177),
	.C1(MK[35]),
	.B2(n188),
	.B1(MK[3]),
	.A2(n205),
	.A1(mkx0[3]));
   OR3B2CHD U227 (
	.O(n504),
	.I1(n267),
	.B2(n269),
	.B1(n268));
   NR3BHD U228 (
	.O(n269),
	.I3(n272),
	.I2(n271),
	.I1(n270));
   OAI22CHD U229 (
	.O(n272),
	.B2(n274),
	.B1(n5),
	.A2(n273),
	.A1(n6));
   OAI222BHD U230 (
	.O(n271),
	.C2(n277),
	.C1(n2),
	.B2(n276),
	.B1(n121),
	.A2(n275),
	.A1(n3));
   AO2222BHD U231 (
	.O(n270),
	.D2(n143),
	.D1(MK[114]),
	.C2(n55),
	.C1(MK[18]),
	.B2(n178),
	.B1(MK[50]),
	.A2(n27),
	.A1(MK[90]));
   OA2222CHD U232 (
	.O(n268),
	.D2(n281),
	.D1(n120),
	.C2(n280),
	.C1(n4),
	.B2(n279),
	.B1(n118),
	.A2(n278),
	.A1(n126));
   AO2222BHD U233 (
	.O(n267),
	.D2(n206),
	.D1(MK[66]),
	.C2(n177),
	.C1(MK[34]),
	.B2(n188),
	.B1(MK[2]),
	.A2(n205),
	.A1(mkx0[2]));
   OR3B2CHD U234 (
	.O(n503),
	.I1(n282),
	.B2(n284),
	.B1(n283));
   NR3BHD U235 (
	.O(n284),
	.I3(n287),
	.I2(n286),
	.I1(n285));
   OAI22CHD U236 (
	.O(n287),
	.B2(n289),
	.B1(n5),
	.A2(n288),
	.A1(n6));
   OAI222BHD U237 (
	.O(n286),
	.C2(n292),
	.C1(n2),
	.B2(n291),
	.B1(n121),
	.A2(n290),
	.A1(n3));
   AO2222BHD U238 (
	.O(n285),
	.D2(n143),
	.D1(MK[113]),
	.C2(n55),
	.C1(MK[17]),
	.B2(n178),
	.B1(MK[49]),
	.A2(n27),
	.A1(MK[89]));
   OA2222CHD U239 (
	.O(n283),
	.D2(n296),
	.D1(n120),
	.C2(n295),
	.C1(n4),
	.B2(n294),
	.B1(n118),
	.A2(n293),
	.A1(n126));
   AO2222BHD U240 (
	.O(n282),
	.D2(n206),
	.D1(MK[65]),
	.C2(n177),
	.C1(MK[33]),
	.B2(n188),
	.B1(MK[1]),
	.A2(n205),
	.A1(mkx0[1]));
   OR3B2CHD U241 (
	.O(n502),
	.I1(n297),
	.B2(n299),
	.B1(n298));
   NR3BHD U242 (
	.O(n299),
	.I3(n302),
	.I2(n301),
	.I1(n300));
   OAI22CHD U243 (
	.O(n302),
	.B2(n304),
	.B1(n5),
	.A2(n303),
	.A1(n6));
   OAI222BHD U244 (
	.O(n301),
	.C2(n307),
	.C1(n2),
	.B2(n306),
	.B1(n121),
	.A2(n305),
	.A1(n3));
   AO2222BHD U245 (
	.O(n300),
	.D2(n143),
	.D1(MK[112]),
	.C2(n55),
	.C1(MK[16]),
	.B2(n178),
	.B1(MK[48]),
	.A2(n27),
	.A1(MK[88]));
   OA2222CHD U246 (
	.O(n298),
	.D2(n311),
	.D1(n120),
	.C2(n310),
	.C1(n4),
	.B2(n309),
	.B1(n118),
	.A2(n308),
	.A1(n126));
   AO2222BHD U247 (
	.O(n297),
	.D2(n206),
	.D1(MK[64]),
	.C2(n177),
	.C1(MK[32]),
	.B2(n188),
	.B1(MK[0]),
	.A2(n205),
	.A1(mkx0[0]));
   OR3B2CHD U248 (
	.O(n501),
	.I1(n312),
	.B2(n314),
	.B1(n313));
   NR3BHD U249 (
	.O(n314),
	.I3(n317),
	.I2(n316),
	.I1(n315));
   OAI22CHD U250 (
	.O(n317),
	.B2(n198),
	.B1(n5),
	.A2(n318),
	.A1(n6));
   OAI222BHD U251 (
	.O(n316),
	.C2(n321),
	.C1(n2),
	.B2(n320),
	.B1(n121),
	.A2(n319),
	.A1(n3));
   AO2222BHD U252 (
	.O(n315),
	.D2(n143),
	.D1(MK[127]),
	.C2(n55),
	.C1(MK[31]),
	.B2(n178),
	.B1(MK[63]),
	.A2(n27),
	.A1(MK[103]));
   OA2222CHD U253 (
	.O(n313),
	.D2(n324),
	.D1(n120),
	.C2(n323),
	.C1(n4),
	.B2(n322),
	.B1(n118),
	.A2(n196),
	.A1(n126));
   AO2222BHD U254 (
	.O(n312),
	.D2(n206),
	.D1(MK[79]),
	.C2(n177),
	.C1(MK[47]),
	.B2(n188),
	.B1(MK[15]),
	.A2(n205),
	.A1(mkx1[7]));
   OR3B2CHD U255 (
	.O(n500),
	.I1(n325),
	.B2(n327),
	.B1(n326));
   NR3BHD U256 (
	.O(n327),
	.I3(n330),
	.I2(n329),
	.I1(n328));
   OAI22CHD U257 (
	.O(n330),
	.B2(n215),
	.B1(n5),
	.A2(n331),
	.A1(n6));
   OAI222BHD U258 (
	.O(n329),
	.C2(n334),
	.C1(n2),
	.B2(n333),
	.B1(n121),
	.A2(n332),
	.A1(n3));
   AO2222BHD U259 (
	.O(n328),
	.D2(n143),
	.D1(MK[126]),
	.C2(n55),
	.C1(MK[30]),
	.B2(n178),
	.B1(MK[62]),
	.A2(n27),
	.A1(MK[102]));
   OA2222CHD U260 (
	.O(n326),
	.D2(n337),
	.D1(n120),
	.C2(n336),
	.C1(n4),
	.B2(n335),
	.B1(n118),
	.A2(n213),
	.A1(n126));
   AO2222BHD U261 (
	.O(n325),
	.D2(n206),
	.D1(MK[78]),
	.C2(n177),
	.C1(MK[46]),
	.B2(n188),
	.B1(MK[14]),
	.A2(n205),
	.A1(mkx1[6]));
   OR3B2CHD U262 (
	.O(n499),
	.I1(n338),
	.B2(n340),
	.B1(n339));
   NR3BHD U263 (
	.O(n340),
	.I3(n343),
	.I2(n342),
	.I1(n341));
   OAI22CHD U264 (
	.O(n343),
	.B2(n230),
	.B1(n5),
	.A2(n344),
	.A1(n6));
   OAI222BHD U265 (
	.O(n342),
	.C2(n347),
	.C1(n2),
	.B2(n346),
	.B1(n121),
	.A2(n345),
	.A1(n3));
   AO2222BHD U266 (
	.O(n341),
	.D2(n143),
	.D1(MK[125]),
	.C2(n55),
	.C1(MK[29]),
	.B2(n178),
	.B1(MK[61]),
	.A2(n27),
	.A1(MK[101]));
   OA2222CHD U267 (
	.O(n339),
	.D2(n350),
	.D1(n120),
	.C2(n349),
	.C1(n4),
	.B2(n348),
	.B1(n118),
	.A2(n228),
	.A1(n126));
   AO2222BHD U268 (
	.O(n338),
	.D2(n206),
	.D1(MK[77]),
	.C2(n177),
	.C1(MK[45]),
	.B2(n188),
	.B1(MK[13]),
	.A2(n205),
	.A1(mkx1[5]));
   OR3B2CHD U269 (
	.O(n498),
	.I1(n351),
	.B2(n353),
	.B1(n352));
   NR3BHD U270 (
	.O(n353),
	.I3(n356),
	.I2(n355),
	.I1(n354));
   OAI22CHD U271 (
	.O(n356),
	.B2(n245),
	.B1(n5),
	.A2(n357),
	.A1(n6));
   OAI222BHD U272 (
	.O(n355),
	.C2(n360),
	.C1(n2),
	.B2(n359),
	.B1(n121),
	.A2(n358),
	.A1(n3));
   AO2222BHD U273 (
	.O(n354),
	.D2(n143),
	.D1(MK[124]),
	.C2(n55),
	.C1(MK[28]),
	.B2(n178),
	.B1(MK[60]),
	.A2(n27),
	.A1(MK[100]));
   OA2222CHD U274 (
	.O(n352),
	.D2(n363),
	.D1(n120),
	.C2(n362),
	.C1(n4),
	.B2(n361),
	.B1(n118),
	.A2(n243),
	.A1(n126));
   AO2222BHD U275 (
	.O(n351),
	.D2(n206),
	.D1(MK[76]),
	.C2(n177),
	.C1(MK[44]),
	.B2(n188),
	.B1(MK[12]),
	.A2(n205),
	.A1(mkx1[4]));
   OR3B2CHD U276 (
	.O(n497),
	.I1(n364),
	.B2(n366),
	.B1(n365));
   NR3BHD U277 (
	.O(n366),
	.I3(n369),
	.I2(n368),
	.I1(n367));
   OAI22CHD U278 (
	.O(n369),
	.B2(n260),
	.B1(n5),
	.A2(n370),
	.A1(n6));
   OAI222BHD U279 (
	.O(n368),
	.C2(n373),
	.C1(n2),
	.B2(n372),
	.B1(n121),
	.A2(n371),
	.A1(n3));
   AO2222BHD U280 (
	.O(n367),
	.D2(n143),
	.D1(MK[123]),
	.C2(n55),
	.C1(MK[27]),
	.B2(n178),
	.B1(MK[59]),
	.A2(n27),
	.A1(MK[99]));
   OA2222CHD U281 (
	.O(n365),
	.D2(n376),
	.D1(n120),
	.C2(n375),
	.C1(n4),
	.B2(n374),
	.B1(n118),
	.A2(n258),
	.A1(n126));
   AO2222BHD U282 (
	.O(n364),
	.D2(n206),
	.D1(MK[75]),
	.C2(n177),
	.C1(MK[43]),
	.B2(n188),
	.B1(MK[11]),
	.A2(n205),
	.A1(mkx1[3]));
   OR3B2CHD U283 (
	.O(n496),
	.I1(n377),
	.B2(n379),
	.B1(n378));
   NR3BHD U284 (
	.O(n379),
	.I3(n382),
	.I2(n381),
	.I1(n380));
   OAI22CHD U285 (
	.O(n382),
	.B2(n275),
	.B1(n5),
	.A2(n383),
	.A1(n6));
   OAI222BHD U286 (
	.O(n381),
	.C2(n386),
	.C1(n2),
	.B2(n385),
	.B1(n121),
	.A2(n384),
	.A1(n3));
   AO2222BHD U287 (
	.O(n380),
	.D2(n143),
	.D1(MK[122]),
	.C2(n55),
	.C1(MK[26]),
	.B2(n178),
	.B1(MK[58]),
	.A2(n27),
	.A1(MK[98]));
   OA2222CHD U288 (
	.O(n378),
	.D2(n389),
	.D1(n120),
	.C2(n388),
	.C1(n4),
	.B2(n387),
	.B1(n118),
	.A2(n273),
	.A1(n126));
   AO2222BHD U289 (
	.O(n377),
	.D2(n206),
	.D1(MK[74]),
	.C2(n177),
	.C1(MK[42]),
	.B2(n188),
	.B1(MK[10]),
	.A2(n205),
	.A1(mkx1[2]));
   OR3B2CHD U290 (
	.O(n495),
	.I1(n390),
	.B2(n392),
	.B1(n391));
   NR3BHD U291 (
	.O(n392),
	.I3(n395),
	.I2(n394),
	.I1(n393));
   OAI22CHD U292 (
	.O(n395),
	.B2(n290),
	.B1(n5),
	.A2(n396),
	.A1(n6));
   OAI222BHD U293 (
	.O(n394),
	.C2(n399),
	.C1(n2),
	.B2(n398),
	.B1(n121),
	.A2(n397),
	.A1(n3));
   AO2222BHD U294 (
	.O(n393),
	.D2(n143),
	.D1(MK[121]),
	.C2(n55),
	.C1(MK[25]),
	.B2(n178),
	.B1(MK[57]),
	.A2(n27),
	.A1(MK[97]));
   OA2222CHD U295 (
	.O(n391),
	.D2(n402),
	.D1(n120),
	.C2(n401),
	.C1(n4),
	.B2(n400),
	.B1(n118),
	.A2(n288),
	.A1(n126));
   AO2222BHD U296 (
	.O(n390),
	.D2(n206),
	.D1(MK[73]),
	.C2(n177),
	.C1(MK[41]),
	.B2(n188),
	.B1(MK[9]),
	.A2(n205),
	.A1(mkx1[1]));
   OR3B2CHD U297 (
	.O(n494),
	.I1(n403),
	.B2(n405),
	.B1(n404));
   NR3BHD U298 (
	.O(n405),
	.I3(n408),
	.I2(n407),
	.I1(n406));
   OAI22CHD U299 (
	.O(n408),
	.B2(n305),
	.B1(n5),
	.A2(n409),
	.A1(n6));
   OAI222BHD U300 (
	.O(n407),
	.C2(n412),
	.C1(n2),
	.B2(n411),
	.B1(n121),
	.A2(n410),
	.A1(n3));
   AO2222BHD U301 (
	.O(n406),
	.D2(n143),
	.D1(MK[120]),
	.C2(n55),
	.C1(MK[24]),
	.B2(n178),
	.B1(MK[56]),
	.A2(n27),
	.A1(MK[96]));
   OA2222CHD U302 (
	.O(n404),
	.D2(n415),
	.D1(n120),
	.C2(n414),
	.C1(n4),
	.B2(n413),
	.B1(n118),
	.A2(n303),
	.A1(n126));
   AO2222BHD U303 (
	.O(n403),
	.D2(n206),
	.D1(MK[72]),
	.C2(n177),
	.C1(MK[40]),
	.B2(n188),
	.B1(MK[8]),
	.A2(n205),
	.A1(mkx1[0]));
   OR3B2CHD U304 (
	.O(n493),
	.I1(n416),
	.B2(n418),
	.B1(n417));
   NR3BHD U305 (
	.O(n418),
	.I3(n421),
	.I2(n420),
	.I1(n419));
   OAI22CHD U306 (
	.O(n421),
	.B2(n319),
	.B1(n5),
	.A2(n204),
	.A1(n6));
   INVCHD U307 (
	.O(n319),
	.I(MK[95]));
   OAI222BHD U308 (
	.O(n420),
	.C2(n203),
	.C1(n2),
	.B2(n202),
	.B1(n121),
	.A2(n201),
	.A1(n3));
   INVCHD U309 (
	.O(n203),
	.I(MK[31]));
   INVCHD U310 (
	.O(n202),
	.I(MK[63]));
   AO2222BHD U311 (
	.O(n419),
	.D2(n143),
	.D1(MK[71]),
	.C2(n55),
	.C1(MK[39]),
	.B2(n178),
	.B1(MK[7]),
	.A2(n27),
	.A1(MK[111]));
   OA2222CHD U312 (
	.O(n417),
	.D2(n197),
	.D1(n120),
	.C2(n199),
	.C1(n4),
	.B2(n200),
	.B1(n118),
	.A2(n318),
	.A1(n126));
   INVCHD U313 (
	.O(n197),
	.I(MK[79]));
   INVCHD U314 (
	.O(n199),
	.I(MK[47]));
   INVCHD U315 (
	.O(n200),
	.I(MK[15]));
   INVCHD U316 (
	.O(n318),
	.I(MK[119]));
   AO2222BHD U317 (
	.O(n416),
	.D2(n206),
	.D1(MK[87]),
	.C2(n177),
	.C1(MK[55]),
	.B2(n188),
	.B1(MK[23]),
	.A2(n205),
	.A1(mkx2[7]));
   OR3B2CHD U318 (
	.O(n492),
	.I1(n422),
	.B2(n424),
	.B1(n423));
   NR3BHD U319 (
	.O(n424),
	.I3(n427),
	.I2(n426),
	.I1(n425));
   OAI22CHD U320 (
	.O(n427),
	.B2(n332),
	.B1(n5),
	.A2(n221),
	.A1(n6));
   INVCHD U321 (
	.O(n332),
	.I(MK[94]));
   OAI222BHD U322 (
	.O(n426),
	.C2(n220),
	.C1(n2),
	.B2(n219),
	.B1(n121),
	.A2(n218),
	.A1(n3));
   INVCHD U323 (
	.O(n220),
	.I(MK[30]));
   INVCHD U324 (
	.O(n219),
	.I(MK[62]));
   AO2222BHD U325 (
	.O(n425),
	.D2(n143),
	.D1(MK[70]),
	.C2(n55),
	.C1(MK[38]),
	.B2(n178),
	.B1(MK[6]),
	.A2(n27),
	.A1(MK[110]));
   OA2222CHD U326 (
	.O(n423),
	.D2(n214),
	.D1(n120),
	.C2(n216),
	.C1(n4),
	.B2(n217),
	.B1(n118),
	.A2(n331),
	.A1(n126));
   INVCHD U327 (
	.O(n214),
	.I(MK[78]));
   INVCHD U328 (
	.O(n216),
	.I(MK[46]));
   INVCHD U329 (
	.O(n217),
	.I(MK[14]));
   INVCHD U330 (
	.O(n331),
	.I(MK[118]));
   AO2222BHD U331 (
	.O(n422),
	.D2(n206),
	.D1(MK[86]),
	.C2(n177),
	.C1(MK[54]),
	.B2(n188),
	.B1(MK[22]),
	.A2(n205),
	.A1(mkx2[6]));
   OR3B2CHD U332 (
	.O(n491),
	.I1(n428),
	.B2(n430),
	.B1(n429));
   NR3BHD U333 (
	.O(n430),
	.I3(n433),
	.I2(n432),
	.I1(n431));
   OAI22CHD U334 (
	.O(n433),
	.B2(n345),
	.B1(n5),
	.A2(n236),
	.A1(n6));
   INVCHD U335 (
	.O(n345),
	.I(MK[93]));
   OAI222BHD U336 (
	.O(n432),
	.C2(n235),
	.C1(n2),
	.B2(n234),
	.B1(n121),
	.A2(n233),
	.A1(n3));
   INVCHD U337 (
	.O(n235),
	.I(MK[29]));
   INVCHD U338 (
	.O(n234),
	.I(MK[61]));
   AO2222BHD U339 (
	.O(n431),
	.D2(n143),
	.D1(MK[69]),
	.C2(n55),
	.C1(MK[37]),
	.B2(n178),
	.B1(MK[5]),
	.A2(n27),
	.A1(MK[109]));
   OA2222CHD U340 (
	.O(n429),
	.D2(n229),
	.D1(n120),
	.C2(n231),
	.C1(n4),
	.B2(n232),
	.B1(n118),
	.A2(n344),
	.A1(n126));
   INVCHD U341 (
	.O(n229),
	.I(MK[77]));
   INVCHD U342 (
	.O(n231),
	.I(MK[45]));
   INVCHD U343 (
	.O(n232),
	.I(MK[13]));
   INVCHD U344 (
	.O(n344),
	.I(MK[117]));
   AO2222BHD U345 (
	.O(n428),
	.D2(n206),
	.D1(MK[85]),
	.C2(n177),
	.C1(MK[53]),
	.B2(n188),
	.B1(MK[21]),
	.A2(n205),
	.A1(mkx2[5]));
   OR3B2CHD U346 (
	.O(n490),
	.I1(n434),
	.B2(n436),
	.B1(n435));
   NR3BHD U347 (
	.O(n436),
	.I3(n439),
	.I2(n438),
	.I1(n437));
   OAI22CHD U348 (
	.O(n439),
	.B2(n358),
	.B1(n5),
	.A2(n251),
	.A1(n6));
   INVCHD U349 (
	.O(n358),
	.I(MK[92]));
   OAI222BHD U350 (
	.O(n438),
	.C2(n250),
	.C1(n2),
	.B2(n249),
	.B1(n121),
	.A2(n248),
	.A1(n3));
   INVCHD U351 (
	.O(n250),
	.I(MK[28]));
   INVCHD U352 (
	.O(n249),
	.I(MK[60]));
   AO2222BHD U353 (
	.O(n437),
	.D2(n143),
	.D1(MK[68]),
	.C2(n55),
	.C1(MK[36]),
	.B2(n178),
	.B1(MK[4]),
	.A2(n27),
	.A1(MK[108]));
   OA2222CHD U354 (
	.O(n435),
	.D2(n244),
	.D1(n120),
	.C2(n246),
	.C1(n4),
	.B2(n247),
	.B1(n118),
	.A2(n357),
	.A1(n126));
   INVCHD U355 (
	.O(n244),
	.I(MK[76]));
   INVCHD U356 (
	.O(n246),
	.I(MK[44]));
   INVCHD U357 (
	.O(n247),
	.I(MK[12]));
   INVCHD U358 (
	.O(n357),
	.I(MK[116]));
   AO2222BHD U359 (
	.O(n434),
	.D2(n206),
	.D1(MK[84]),
	.C2(n177),
	.C1(MK[52]),
	.B2(n188),
	.B1(MK[20]),
	.A2(n205),
	.A1(mkx2[4]));
   OR3B2CHD U360 (
	.O(n489),
	.I1(n440),
	.B2(n442),
	.B1(n441));
   NR3BHD U361 (
	.O(n442),
	.I3(n445),
	.I2(n444),
	.I1(n443));
   OAI22CHD U362 (
	.O(n445),
	.B2(n371),
	.B1(n5),
	.A2(n266),
	.A1(n6));
   INVCHD U363 (
	.O(n371),
	.I(MK[91]));
   OAI222BHD U364 (
	.O(n444),
	.C2(n265),
	.C1(n2),
	.B2(n264),
	.B1(n121),
	.A2(n263),
	.A1(n3));
   INVCHD U365 (
	.O(n265),
	.I(MK[27]));
   INVCHD U366 (
	.O(n264),
	.I(MK[59]));
   AO2222BHD U367 (
	.O(n443),
	.D2(n143),
	.D1(MK[67]),
	.C2(n55),
	.C1(MK[35]),
	.B2(n178),
	.B1(MK[3]),
	.A2(n27),
	.A1(MK[107]));
   OA2222CHD U368 (
	.O(n441),
	.D2(n259),
	.D1(n120),
	.C2(n261),
	.C1(n4),
	.B2(n262),
	.B1(n118),
	.A2(n370),
	.A1(n126));
   INVCHD U369 (
	.O(n259),
	.I(MK[75]));
   INVCHD U370 (
	.O(n261),
	.I(MK[43]));
   INVCHD U371 (
	.O(n262),
	.I(MK[11]));
   INVCHD U372 (
	.O(n370),
	.I(MK[115]));
   AO2222BHD U373 (
	.O(n440),
	.D2(n206),
	.D1(MK[83]),
	.C2(n177),
	.C1(MK[51]),
	.B2(n188),
	.B1(MK[19]),
	.A2(n205),
	.A1(mkx2[3]));
   OR3B2CHD U374 (
	.O(n488),
	.I1(n446),
	.B2(n448),
	.B1(n447));
   NR3BHD U375 (
	.O(n448),
	.I3(n451),
	.I2(n450),
	.I1(n449));
   OAI22CHD U376 (
	.O(n451),
	.B2(n384),
	.B1(n5),
	.A2(n281),
	.A1(n6));
   INVCHD U377 (
	.O(n384),
	.I(MK[90]));
   OAI222BHD U378 (
	.O(n450),
	.C2(n280),
	.C1(n2),
	.B2(n279),
	.B1(n121),
	.A2(n278),
	.A1(n3));
   INVCHD U379 (
	.O(n280),
	.I(MK[26]));
   INVCHD U380 (
	.O(n279),
	.I(MK[58]));
   AO2222BHD U381 (
	.O(n449),
	.D2(n143),
	.D1(MK[66]),
	.C2(n55),
	.C1(MK[34]),
	.B2(n178),
	.B1(MK[2]),
	.A2(n27),
	.A1(MK[106]));
   OA2222CHD U382 (
	.O(n447),
	.D2(n274),
	.D1(n120),
	.C2(n276),
	.C1(n4),
	.B2(n277),
	.B1(n118),
	.A2(n383),
	.A1(n126));
   INVCHD U383 (
	.O(n274),
	.I(MK[74]));
   INVCHD U384 (
	.O(n276),
	.I(MK[42]));
   INVCHD U385 (
	.O(n277),
	.I(MK[10]));
   INVCHD U386 (
	.O(n383),
	.I(MK[114]));
   AO2222BHD U387 (
	.O(n446),
	.D2(n206),
	.D1(MK[82]),
	.C2(n177),
	.C1(MK[50]),
	.B2(n188),
	.B1(MK[18]),
	.A2(n205),
	.A1(mkx2[2]));
   OR3B2CHD U388 (
	.O(n487),
	.I1(n452),
	.B2(n454),
	.B1(n453));
   NR3BHD U389 (
	.O(n454),
	.I3(n457),
	.I2(n456),
	.I1(n455));
   OAI22CHD U390 (
	.O(n457),
	.B2(n397),
	.B1(n5),
	.A2(n296),
	.A1(n6));
   INVCHD U391 (
	.O(n397),
	.I(MK[89]));
   OAI222BHD U392 (
	.O(n456),
	.C2(n295),
	.C1(n2),
	.B2(n294),
	.B1(n121),
	.A2(n293),
	.A1(n3));
   INVCHD U393 (
	.O(n295),
	.I(MK[25]));
   INVCHD U394 (
	.O(n294),
	.I(MK[57]));
   AO2222BHD U395 (
	.O(n455),
	.D2(n143),
	.D1(MK[65]),
	.C2(n55),
	.C1(MK[33]),
	.B2(n178),
	.B1(MK[1]),
	.A2(n27),
	.A1(MK[105]));
   OA2222CHD U396 (
	.O(n453),
	.D2(n289),
	.D1(n120),
	.C2(n291),
	.C1(n4),
	.B2(n292),
	.B1(n118),
	.A2(n396),
	.A1(n126));
   INVCHD U397 (
	.O(n289),
	.I(MK[73]));
   INVCHD U398 (
	.O(n291),
	.I(MK[41]));
   INVCHD U399 (
	.O(n292),
	.I(MK[9]));
   INVCHD U400 (
	.O(n396),
	.I(MK[113]));
   AO2222BHD U401 (
	.O(n452),
	.D2(n206),
	.D1(MK[81]),
	.C2(n177),
	.C1(MK[49]),
	.B2(n188),
	.B1(MK[17]),
	.A2(n205),
	.A1(mkx2[1]));
   OR3B2CHD U402 (
	.O(n486),
	.I1(n458),
	.B2(n460),
	.B1(n459));
   NR3BHD U403 (
	.O(n460),
	.I3(n463),
	.I2(n462),
	.I1(n461));
   OAI22CHD U404 (
	.O(n463),
	.B2(n410),
	.B1(n5),
	.A2(n311),
	.A1(n6));
   INVCHD U405 (
	.O(n410),
	.I(MK[88]));
   OAI222BHD U406 (
	.O(n462),
	.C2(n310),
	.C1(n2),
	.B2(n309),
	.B1(n121),
	.A2(n308),
	.A1(n3));
   INVCHD U407 (
	.O(n310),
	.I(MK[24]));
   INVCHD U408 (
	.O(n309),
	.I(MK[56]));
   AO2222BHD U409 (
	.O(n461),
	.D2(n143),
	.D1(MK[64]),
	.C2(n55),
	.C1(MK[32]),
	.B2(n178),
	.B1(MK[0]),
	.A2(n27),
	.A1(MK[104]));
   OA2222CHD U410 (
	.O(n459),
	.D2(n304),
	.D1(n120),
	.C2(n306),
	.C1(n4),
	.B2(n307),
	.B1(n118),
	.A2(n409),
	.A1(n126));
   INVCHD U411 (
	.O(n304),
	.I(MK[72]));
   INVCHD U412 (
	.O(n306),
	.I(MK[40]));
   INVCHD U413 (
	.O(n307),
	.I(MK[8]));
   INVCHD U414 (
	.O(n409),
	.I(MK[112]));
   AO2222BHD U415 (
	.O(n458),
	.D2(n206),
	.D1(MK[80]),
	.C2(n177),
	.C1(MK[48]),
	.B2(n188),
	.B1(MK[16]),
	.A2(n205),
	.A1(mkx2[0]));
   OR3B2CHD U416 (
	.O(n485),
	.I1(n464),
	.B2(n466),
	.B1(n465));
   NR3BHD U417 (
	.O(n466),
	.I3(n469),
	.I2(n468),
	.I1(n467));
   OAI22CHD U418 (
	.O(n469),
	.B2(n201),
	.B1(n5),
	.A2(n324),
	.A1(n6));
   INVCHD U419 (
	.O(n201),
	.I(MK[103]));
   INVCHD U420 (
	.O(n324),
	.I(MK[71]));
   OAI222BHD U421 (
	.O(n468),
	.C2(n323),
	.C1(n2),
	.B2(n322),
	.B1(n121),
	.A2(n196),
	.A1(n3));
   INVCHD U422 (
	.O(n323),
	.I(MK[39]));
   INVCHD U423 (
	.O(n322),
	.I(MK[7]));
   INVCHD U424 (
	.O(n196),
	.I(MK[111]));
   AO2222BHD U425 (
	.O(n467),
	.D2(n143),
	.D1(MK[79]),
	.C2(n55),
	.C1(MK[47]),
	.B2(n178),
	.B1(MK[15]),
	.A2(n27),
	.A1(MK[119]));
   OA2222CHD U426 (
	.O(n465),
	.D2(n198),
	.D1(n120),
	.C2(n320),
	.C1(n4),
	.B2(n321),
	.B1(n118),
	.A2(n204),
	.A1(n126));
   INVCHD U427 (
	.O(n198),
	.I(MK[87]));
   INVCHD U428 (
	.O(n320),
	.I(MK[55]));
   INVCHD U429 (
	.O(n321),
	.I(MK[23]));
   INVCHD U430 (
	.O(n204),
	.I(MK[127]));
   AO2222BHD U431 (
	.O(n464),
	.D2(n206),
	.D1(MK[95]),
	.C2(n177),
	.C1(MK[63]),
	.B2(n188),
	.B1(MK[31]),
	.A2(n205),
	.A1(mkx3[7]));
   OR3B2CHD U432 (
	.O(n484),
	.I1(n470),
	.B2(n472),
	.B1(n471));
   NR3BHD U433 (
	.O(n472),
	.I3(n475),
	.I2(n474),
	.I1(n473));
   OAI22CHD U434 (
	.O(n475),
	.B2(n218),
	.B1(n5),
	.A2(n337),
	.A1(n6));
   INVCHD U435 (
	.O(n218),
	.I(MK[102]));
   INVCHD U436 (
	.O(n337),
	.I(MK[70]));
   OAI222BHD U437 (
	.O(n474),
	.C2(n336),
	.C1(n2),
	.B2(n335),
	.B1(n121),
	.A2(n213),
	.A1(n3));
   INVCHD U438 (
	.O(n336),
	.I(MK[38]));
   INVCHD U439 (
	.O(n335),
	.I(MK[6]));
   INVCHD U440 (
	.O(n213),
	.I(MK[110]));
   AO2222BHD U441 (
	.O(n473),
	.D2(n143),
	.D1(MK[78]),
	.C2(n55),
	.C1(MK[46]),
	.B2(n178),
	.B1(MK[14]),
	.A2(n27),
	.A1(MK[118]));
   OA2222CHD U442 (
	.O(n471),
	.D2(n215),
	.D1(n120),
	.C2(n333),
	.C1(n4),
	.B2(n334),
	.B1(n118),
	.A2(n221),
	.A1(n126));
   INVCHD U443 (
	.O(n215),
	.I(MK[86]));
   INVCHD U444 (
	.O(n333),
	.I(MK[54]));
   INVCHD U445 (
	.O(n334),
	.I(MK[22]));
   INVCHD U446 (
	.O(n221),
	.I(MK[126]));
   AO2222BHD U447 (
	.O(n470),
	.D2(n206),
	.D1(MK[94]),
	.C2(n177),
	.C1(MK[62]),
	.B2(n188),
	.B1(MK[30]),
	.A2(n205),
	.A1(mkx3[6]));
   OR3B2CHD U448 (
	.O(n483),
	.I1(n476),
	.B2(n544),
	.B1(n477));
   NR3BHD U449 (
	.O(n544),
	.I3(n547),
	.I2(n546),
	.I1(n545));
   OAI22CHD U450 (
	.O(n547),
	.B2(n233),
	.B1(n5),
	.A2(n350),
	.A1(n6));
   INVCHD U451 (
	.O(n233),
	.I(MK[101]));
   INVCHD U452 (
	.O(n350),
	.I(MK[69]));
   OAI222BHD U453 (
	.O(n546),
	.C2(n349),
	.C1(n2),
	.B2(n348),
	.B1(n121),
	.A2(n228),
	.A1(n3));
   INVCHD U454 (
	.O(n349),
	.I(MK[37]));
   INVCHD U455 (
	.O(n348),
	.I(MK[5]));
   INVCHD U456 (
	.O(n228),
	.I(MK[109]));
   AO2222BHD U457 (
	.O(n545),
	.D2(n143),
	.D1(MK[77]),
	.C2(n55),
	.C1(MK[45]),
	.B2(n178),
	.B1(MK[13]),
	.A2(n27),
	.A1(MK[117]));
   OA2222CHD U458 (
	.O(n477),
	.D2(n230),
	.D1(n120),
	.C2(n346),
	.C1(n4),
	.B2(n347),
	.B1(n118),
	.A2(n236),
	.A1(n126));
   INVCHD U459 (
	.O(n230),
	.I(MK[85]));
   INVCHD U460 (
	.O(n346),
	.I(MK[53]));
   INVCHD U461 (
	.O(n347),
	.I(MK[21]));
   INVCHD U462 (
	.O(n236),
	.I(MK[125]));
   AO2222BHD U463 (
	.O(n476),
	.D2(n206),
	.D1(MK[93]),
	.C2(n177),
	.C1(MK[61]),
	.B2(n188),
	.B1(MK[29]),
	.A2(n205),
	.A1(mkx3[5]));
   OR3B2CHD U464 (
	.O(n482),
	.I1(n548),
	.B2(n550),
	.B1(n549));
   NR3BHD U465 (
	.O(n550),
	.I3(n553),
	.I2(n552),
	.I1(n551));
   OAI22CHD U466 (
	.O(n553),
	.B2(n248),
	.B1(n5),
	.A2(n363),
	.A1(n6));
   INVCHD U467 (
	.O(n248),
	.I(MK[100]));
   INVCHD U468 (
	.O(n363),
	.I(MK[68]));
   OAI222BHD U469 (
	.O(n552),
	.C2(n362),
	.C1(n2),
	.B2(n361),
	.B1(n121),
	.A2(n243),
	.A1(n3));
   INVCHD U470 (
	.O(n362),
	.I(MK[36]));
   INVCHD U471 (
	.O(n361),
	.I(MK[4]));
   INVCHD U472 (
	.O(n243),
	.I(MK[108]));
   AO2222BHD U473 (
	.O(n551),
	.D2(n143),
	.D1(MK[76]),
	.C2(n55),
	.C1(MK[44]),
	.B2(n178),
	.B1(MK[12]),
	.A2(n27),
	.A1(MK[116]));
   OA2222CHD U474 (
	.O(n549),
	.D2(n245),
	.D1(n120),
	.C2(n359),
	.C1(n4),
	.B2(n360),
	.B1(n118),
	.A2(n251),
	.A1(n126));
   INVCHD U475 (
	.O(n245),
	.I(MK[84]));
   INVCHD U476 (
	.O(n359),
	.I(MK[52]));
   INVCHD U477 (
	.O(n360),
	.I(MK[20]));
   INVCHD U478 (
	.O(n251),
	.I(MK[124]));
   AO2222BHD U479 (
	.O(n548),
	.D2(n206),
	.D1(MK[92]),
	.C2(n177),
	.C1(MK[60]),
	.B2(n188),
	.B1(MK[28]),
	.A2(n205),
	.A1(mkx3[4]));
   OR3B2CHD U480 (
	.O(n481),
	.I1(n554),
	.B2(n556),
	.B1(n555));
   NR3BHD U481 (
	.O(n556),
	.I3(n559),
	.I2(n558),
	.I1(n557));
   OAI22CHD U482 (
	.O(n559),
	.B2(n263),
	.B1(n5),
	.A2(n376),
	.A1(n6));
   INVCHD U483 (
	.O(n263),
	.I(MK[99]));
   INVCHD U484 (
	.O(n376),
	.I(MK[67]));
   OAI222BHD U485 (
	.O(n558),
	.C2(n375),
	.C1(n2),
	.B2(n374),
	.B1(n121),
	.A2(n258),
	.A1(n3));
   INVCHD U486 (
	.O(n375),
	.I(MK[35]));
   INVCHD U487 (
	.O(n374),
	.I(MK[3]));
   INVCHD U488 (
	.O(n258),
	.I(MK[107]));
   AO2222BHD U489 (
	.O(n557),
	.D2(n143),
	.D1(MK[75]),
	.C2(n55),
	.C1(MK[43]),
	.B2(n178),
	.B1(MK[11]),
	.A2(n27),
	.A1(MK[115]));
   OA2222CHD U490 (
	.O(n555),
	.D2(n260),
	.D1(n120),
	.C2(n372),
	.C1(n4),
	.B2(n373),
	.B1(n118),
	.A2(n266),
	.A1(n126));
   INVCHD U491 (
	.O(n260),
	.I(MK[83]));
   INVCHD U492 (
	.O(n372),
	.I(MK[51]));
   INVCHD U493 (
	.O(n373),
	.I(MK[19]));
   INVCHD U494 (
	.O(n266),
	.I(MK[123]));
   AO2222BHD U495 (
	.O(n554),
	.D2(n206),
	.D1(MK[91]),
	.C2(n177),
	.C1(MK[59]),
	.B2(n188),
	.B1(MK[27]),
	.A2(n205),
	.A1(mkx3[3]));
   OR3B2CHD U496 (
	.O(n480),
	.I1(n560),
	.B2(n562),
	.B1(n561));
   NR3BHD U497 (
	.O(n562),
	.I3(n565),
	.I2(n564),
	.I1(n563));
   OAI22CHD U498 (
	.O(n565),
	.B2(n278),
	.B1(n5),
	.A2(n389),
	.A1(n6));
   INVCHD U499 (
	.O(n278),
	.I(MK[98]));
   INVCHD U500 (
	.O(n389),
	.I(MK[66]));
   OAI222BHD U501 (
	.O(n564),
	.C2(n388),
	.C1(n2),
	.B2(n387),
	.B1(n121),
	.A2(n273),
	.A1(n3));
   INVCHD U502 (
	.O(n388),
	.I(MK[34]));
   INVCHD U503 (
	.O(n387),
	.I(MK[2]));
   INVCHD U504 (
	.O(n273),
	.I(MK[106]));
   AO2222BHD U505 (
	.O(n563),
	.D2(n143),
	.D1(MK[74]),
	.C2(n55),
	.C1(MK[42]),
	.B2(n178),
	.B1(MK[10]),
	.A2(n27),
	.A1(MK[114]));
   OA2222CHD U506 (
	.O(n561),
	.D2(n275),
	.D1(n120),
	.C2(n385),
	.C1(n4),
	.B2(n386),
	.B1(n118),
	.A2(n281),
	.A1(n126));
   INVCHD U507 (
	.O(n275),
	.I(MK[82]));
   INVCHD U508 (
	.O(n385),
	.I(MK[50]));
   INVCHD U509 (
	.O(n386),
	.I(MK[18]));
   INVCHD U510 (
	.O(n281),
	.I(MK[122]));
   AO2222BHD U511 (
	.O(n560),
	.D2(n206),
	.D1(MK[90]),
	.C2(n177),
	.C1(MK[58]),
	.B2(n188),
	.B1(MK[26]),
	.A2(n205),
	.A1(mkx3[2]));
   OR3B2CHD U512 (
	.O(n479),
	.I1(n566),
	.B2(n568),
	.B1(n567));
   NR3BHD U513 (
	.O(n568),
	.I3(n571),
	.I2(n570),
	.I1(n569));
   OAI22CHD U514 (
	.O(n571),
	.B2(n293),
	.B1(n5),
	.A2(n402),
	.A1(n6));
   INVCHD U515 (
	.O(n293),
	.I(MK[97]));
   INVCHD U516 (
	.O(n402),
	.I(MK[65]));
   OAI222BHD U517 (
	.O(n570),
	.C2(n401),
	.C1(n2),
	.B2(n400),
	.B1(n121),
	.A2(n288),
	.A1(n3));
   INVCHD U518 (
	.O(n401),
	.I(MK[33]));
   INVCHD U519 (
	.O(n400),
	.I(MK[1]));
   INVCHD U520 (
	.O(n288),
	.I(MK[105]));
   AO2222BHD U521 (
	.O(n569),
	.D2(n143),
	.D1(MK[73]),
	.C2(n55),
	.C1(MK[41]),
	.B2(n178),
	.B1(MK[9]),
	.A2(n27),
	.A1(MK[113]));
   OA2222CHD U522 (
	.O(n567),
	.D2(n290),
	.D1(n120),
	.C2(n398),
	.C1(n4),
	.B2(n399),
	.B1(n118),
	.A2(n296),
	.A1(n126));
   INVCHD U523 (
	.O(n290),
	.I(MK[81]));
   INVCHD U524 (
	.O(n398),
	.I(MK[49]));
   INVCHD U525 (
	.O(n399),
	.I(MK[17]));
   INVCHD U526 (
	.O(n296),
	.I(MK[121]));
   AO2222BHD U527 (
	.O(n566),
	.D2(n206),
	.D1(MK[89]),
	.C2(n177),
	.C1(MK[57]),
	.B2(n188),
	.B1(MK[25]),
	.A2(n205),
	.A1(mkx3[1]));
   OR3B2CHD U528 (
	.O(n478),
	.I1(n572),
	.B2(n574),
	.B1(n573));
   NR3BHD U529 (
	.O(n574),
	.I3(n577),
	.I2(n576),
	.I1(n575));
   OAI22CHD U530 (
	.O(n577),
	.B2(n308),
	.B1(n5),
	.A2(n415),
	.A1(n6));
   INVCHD U531 (
	.O(n308),
	.I(MK[96]));
   NR2BHD U532 (
	.O(n140),
	.I2(n92),
	.I1(n578));
   INVCHD U533 (
	.O(n415),
	.I(MK[64]));
   INVCHD U534 (
	.O(n158),
	.I(n187));
   OAI222BHD U535 (
	.O(n576),
	.C2(n414),
	.C1(n2),
	.B2(n413),
	.B1(n121),
	.A2(n303),
	.A1(n3));
   INVCHD U536 (
	.O(n414),
	.I(MK[32]));
   NR2BHD U537 (
	.O(n115),
	.I2(n144),
	.I1(n148));
   INVCHD U538 (
	.O(n413),
	.I(MK[0]));
   OAI12CHD U539 (
	.O(n113),
	.B2(n149),
	.B1(n148),
	.A1(n173));
   ND2CHD U540 (
	.O(n173),
	.I2(n142),
	.I1(n162));
   NR3BHD U541 (
	.O(n162),
	.I3(n581),
	.I2(n580),
	.I1(n579));
   INVCHD U542 (
	.O(n303),
	.I(MK[104]));
   NR2BHD U543 (
	.O(n153),
	.I2(n93),
	.I1(n148));
   AO2222BHD U544 (
	.O(n575),
	.D2(n143),
	.D1(MK[72]),
	.C2(n55),
	.C1(MK[40]),
	.B2(n178),
	.B1(MK[8]),
	.A2(n27),
	.A1(MK[112]));
   OAI12CHD U545 (
	.O(n143),
	.B2(n148),
	.B1(n578),
	.A1(n174));
   INVCHD U546 (
	.O(n174),
	.I(n164));
   NR2BHD U547 (
	.O(n164),
	.I2(n144),
	.I1(n109));
   INVCHD U548 (
	.O(n148),
	.I(n123));
   NR3BHD U549 (
	.O(n123),
	.I3(n581),
	.I2(i_round[0]),
	.I1(n579));
   OAI22CHD U550 (
	.O(n189),
	.B2(n109),
	.B1(n578),
	.A2(n145),
	.A1(n144));
   OAI22CHD U551 (
	.O(n178),
	.B2(n109),
	.B1(n93),
	.A2(n145),
	.A1(n149));
   INVCHD U552 (
	.O(n109),
	.I(n582));
   NR3BHD U553 (
	.O(n582),
	.I3(n581),
	.I2(i_round[2]),
	.I1(n580));
   INVCHD U554 (
	.O(n581),
	.I(i_round[3]));
   ND2CHD U555 (
	.O(n106),
	.I2(n141),
	.I1(n186));
   OA2222CHD U556 (
	.O(n573),
	.D2(n305),
	.D1(n120),
	.C2(n411),
	.C1(n4),
	.B2(n412),
	.B1(n118),
	.A2(n311),
	.A1(n126));
   INVCHD U557 (
	.O(n305),
	.I(MK[80]));
   ND2CHD U558 (
	.O(n138),
	.I2(n141),
	.I1(n133));
   ND3CHD U559 (
	.O(n145),
	.I3(i_round[3]),
	.I2(n579),
	.I1(n580));
   INVCHD U560 (
	.O(n411),
	.I(MK[48]));
   AN2CHD U561 (
	.O(n152),
	.I2(n141),
	.I1(n124));
   INVCHD U562 (
	.O(n412),
	.I(MK[16]));
   NR2BHD U563 (
	.O(n159),
	.I2(n156),
	.I1(n149));
   NR3BHD U564 (
	.O(n141),
	.I3(n579),
	.I2(i_round[3]),
	.I1(n580));
   INVCHD U565 (
	.O(n311),
	.I(MK[120]));
   NR2BHD U566 (
	.O(n170),
	.I2(n149),
	.I1(n171));
   AO2222BHD U567 (
	.O(n572),
	.D2(n206),
	.D1(MK[88]),
	.C2(n177),
	.C1(MK[56]),
	.B2(n188),
	.B1(MK[24]),
	.A2(n205),
	.A1(mkx3[0]));
   INVCHD U568 (
	.O(n206),
	.I(n136));
   NR2BHD U569 (
	.O(n136),
	.I2(n166),
	.I1(n116));
   NR2BHD U570 (
	.O(n166),
	.I2(n144),
	.I1(n171));
   INVCHD U571 (
	.O(n144),
	.I(n133));
   NR2BHD U572 (
	.O(n116),
	.I2(n578),
	.I1(n156));
   INVCHD U573 (
	.O(n578),
	.I(n124));
   INVCHD U574 (
	.O(n156),
	.I(n131));
   NR3BHD U575 (
	.O(n131),
	.I3(n579),
	.I2(i_round[3]),
	.I1(i_round[0]));
   INVCHD U576 (
	.O(n579),
	.I(i_round[2]));
   INVCHD U577 (
	.O(n177),
	.I(n134));
   AOI22BHD U578 (
	.O(n134),
	.B2(n167),
	.B1(n124),
	.A2(n133),
	.A1(n132));
   NR3BHD U579 (
	.O(n133),
	.I3(n584),
	.I2(i_round[5]),
	.I1(i_round[4]));
   OAI12CHD U580 (
	.O(n188),
	.B2(n171),
	.B1(n93),
	.A1(n150));
   INVCHD U581 (
	.O(n150),
	.I(n104));
   NR2BHD U582 (
	.O(n104),
	.I2(n92),
	.I1(n149));
   INVCHD U583 (
	.O(n149),
	.I(n186));
   NR2BHD U584 (
	.O(n186),
	.I2(n584),
	.I1(n583));
   INVCHD U585 (
	.O(n584),
	.I(i_round[1]));
   INVCHD U586 (
	.O(n171),
	.I(n167));
   NR3BHD U587 (
	.O(n167),
	.I3(n580),
	.I2(i_round[3]),
	.I1(i_round[2]));
   INVCHD U588 (
	.O(n580),
	.I(i_round[0]));
   INVCHD U589 (
	.O(n93),
	.I(n142));
   NR2BHD U590 (
	.O(n142),
	.I2(i_round[5]),
	.I1(n91));
   INVCHD U591 (
	.O(n91),
	.I(n585));
   OA112CHD U592 (
	.O(n205),
	.C2(i_round[5]),
	.C1(n586),
	.B1(n187),
	.A1(n583));
   ND3CHD U593 (
	.O(n187),
	.I3(i_round[5]),
	.I2(n585),
	.I1(n132));
   NR2BHD U594 (
	.O(n585),
	.I2(i_round[4]),
	.I1(i_round[1]));
   OR2B1CHD U595 (
	.O(n583),
	.I1(i_round[5]),
	.B1(i_round[4]));
   NR2BHD U596 (
	.O(n586),
	.I2(n92),
	.I1(i_round[1]));
   INVCHD U597 (
	.O(n92),
	.I(n132));
   NR3BHD U598 (
	.O(n132),
	.I3(i_round[0]),
	.I2(i_round[3]),
	.I1(i_round[2]));
endmodule

module round_funct_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   INVDHD U1 (
	.O(n6),
	.I(B[2]));
   INVDHD U2 (
	.O(n7),
	.I(B[1]));
   INVDHD U3 (
	.O(n3),
	.I(B[5]));
   INVDHD U4 (
	.O(n8),
	.I(B[0]));
   INVDHD U5 (
	.O(n5),
	.I(B[3]));
   INVDHD U6 (
	.O(n4),
	.I(B[4]));
   INVDHD U7 (
	.O(n2),
	.I(B[6]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_sub_1 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   INVDHD U1 (
	.O(n1),
	.I(B[7]));
   INVDHD U2 (
	.O(n3),
	.I(B[5]));
   INVDHD U3 (
	.O(n5),
	.I(B[3]));
   INVDHD U4 (
	.O(n4),
	.I(B[4]));
   INVDHD U5 (
	.O(n2),
	.I(B[6]));
   INVDHD U6 (
	.O(n7),
	.I(B[1]));
   INVDHD U7 (
	.O(n6),
	.I(B[2]));
   INVDHD U8 (
	.O(n8),
	.I(B[0]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_sub_2 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   INVDHD U1 (
	.O(n6),
	.I(B[2]));
   INVDHD U2 (
	.O(n3),
	.I(B[5]));
   INVDHD U3 (
	.O(n7),
	.I(B[1]));
   INVDHD U4 (
	.O(n5),
	.I(B[3]));
   INVDHD U5 (
	.O(n4),
	.I(B[4]));
   INVDHD U6 (
	.O(n2),
	.I(B[6]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_add_2 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_sub_3 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   INVDHD U1 (
	.O(n6),
	.I(B[2]));
   INVDHD U2 (
	.O(n3),
	.I(B[5]));
   INVDHD U3 (
	.O(n7),
	.I(B[1]));
   INVDHD U4 (
	.O(n5),
	.I(B[3]));
   INVDHD U5 (
	.O(n4),
	.I(B[4]));
   INVDHD U6 (
	.O(n2),
	.I(B[6]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_add_3 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_sub_4 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   INVDHD U1 (
	.O(n6),
	.I(B[2]));
   INVDHD U2 (
	.O(n5),
	.I(B[3]));
   INVDHD U3 (
	.O(n4),
	.I(B[4]));
   INVDHD U4 (
	.O(n3),
	.I(B[5]));
   INVDHD U5 (
	.O(n2),
	.I(B[6]));
   INVDHD U6 (
	.O(n7),
	.I(B[1]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_sub_5 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   INVDHD U1 (
	.O(n6),
	.I(B[2]));
   INVDHD U2 (
	.O(n3),
	.I(B[5]));
   INVDHD U3 (
	.O(n7),
	.I(B[1]));
   INVDHD U4 (
	.O(n5),
	.I(B[3]));
   INVDHD U5 (
	.O(n4),
	.I(B[4]));
   INVDHD U6 (
	.O(n2),
	.I(B[6]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_sub_6 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   INVDHD U1 (
	.O(n5),
	.I(B[3]));
   INVDHD U2 (
	.O(n6),
	.I(B[2]));
   INVDHD U3 (
	.O(n4),
	.I(B[4]));
   INVDHD U4 (
	.O(n3),
	.I(B[5]));
   INVDHD U5 (
	.O(n2),
	.I(B[6]));
   INVDHD U6 (
	.O(n7),
	.I(B[1]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_add_4 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_sub_7 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] DIFF;
   output CO;

   // Internal wires
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [8:0] carry;

   // Module instantiations
   XOR3EHD U2_7 (
	.O(DIFF[7]),
	.I3(carry[7]),
	.I2(n1),
	.I1(A[7]));
   FA1DHD U2_0 (
	.S(DIFF[0]),
	.CO(carry[1]),
	.CI(n9),
	.B(n8),
	.A(A[0]));
   FA1DHD U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n7),
	.A(A[1]));
   FA1DHD U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n2),
	.A(A[6]));
   FA1DHD U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n3),
	.A(A[5]));
   FA1DHD U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n6),
	.A(A[2]));
   FA1DHD U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n5),
	.A(A[3]));
   FA1DHD U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n4),
	.A(A[4]));
   INVDHD U1 (
	.O(n4),
	.I(B[4]));
   INVDHD U2 (
	.O(n5),
	.I(B[3]));
   INVDHD U3 (
	.O(n6),
	.I(B[2]));
   INVDHD U4 (
	.O(n3),
	.I(B[5]));
   INVDHD U5 (
	.O(n2),
	.I(B[6]));
   INVDHD U6 (
	.O(n7),
	.I(B[1]));
   INVDHD U7 (
	.O(n8),
	.I(B[0]));
   INVDHD U8 (
	.O(n1),
	.I(B[7]));
   TIE1DHD U9 (
	.O(n9));
endmodule

module round_funct_DW01_add_5 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_add_6 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_add_7 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_add_8 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct_DW01_add_9 (
	A, 
	B, 
	CI, 
	SUM, 
	CO);
   input [7:0] A;
   input [7:0] B;
   input CI;
   output [7:0] SUM;
   output CO;

   // Internal wires
   wire n1;
   wire [7:1] carry;

   // Module instantiations
   FA1DHD U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]));
   FA1DHD U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]));
   FA1DHD U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]));
   FA1DHD U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]));
   FA1DHD U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]));
   FA1DHD U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(B[1]),
	.A(A[1]));
   FA1DHD U1_0 (
	.S(SUM[0]),
	.CO(carry[1]),
	.CI(n1),
	.B(B[0]),
	.A(A[0]));
   XOR3EHD U1_7 (
	.O(SUM[7]),
	.I3(carry[7]),
	.I2(B[7]),
	.I1(A[7]));
   TIE0DHD U1 (
	.O(n1));
endmodule

module round_funct (
	P, 
	MK, 
	SKx0, 
	SKx1, 
	SKx2, 
	SKx3, 
	clk, 
	reset, 
	ed, 
	WK0_4, 
	WK1_5, 
	WK2_6, 
	WK3_7, 
	C);
   input [63:0] P;
   input [127:0] MK;
   input [7:0] SKx0;
   input [7:0] SKx1;
   input [7:0] SKx2;
   input [7:0] SKx3;
   input clk;
   input reset;
   input ed;
   input [7:0] WK0_4;
   input [7:0] WK1_5;
   input [7:0] WK2_6;
   input [7:0] WK3_7;
   output [63:0] C;

   // Internal wires
   wire N6;
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N23;
   wire N26;
   wire N27;
   wire N28;
   wire N29;
   wire N30;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire N48;
   wire N49;
   wire N50;
   wire N51;
   wire N52;
   wire N53;
   wire N54;
   wire N55;
   wire N56;
   wire N57;
   wire N58;
   wire N75;
   wire N76;
   wire N77;
   wire N78;
   wire N79;
   wire N80;
   wire N81;
   wire N82;
   wire N83;
   wire N84;
   wire N85;
   wire N86;
   wire N87;
   wire N88;
   wire N89;
   wire N90;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N132;
   wire N133;
   wire N134;
   wire N135;
   wire N136;
   wire N137;
   wire N138;
   wire N139;
   wire N140;
   wire N141;
   wire N142;
   wire N143;
   wire N144;
   wire N145;
   wire N146;
   wire N147;
   wire N173;
   wire N174;
   wire N175;
   wire N176;
   wire N177;
   wire N178;
   wire N179;
   wire N180;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire N201;
   wire N202;
   wire N203;
   wire N204;
   wire N255;
   wire N256;
   wire N257;
   wire N258;
   wire N259;
   wire N260;
   wire N261;
   wire N262;
   wire N263;
   wire N264;
   wire N265;
   wire N266;
   wire N267;
   wire N268;
   wire N269;
   wire N270;
   wire N287;
   wire N288;
   wire N289;
   wire N290;
   wire N291;
   wire N292;
   wire N293;
   wire N294;
   wire N295;
   wire N296;
   wire N297;
   wire N298;
   wire N299;
   wire N300;
   wire N301;
   wire N302;
   wire N389;
   wire N390;
   wire N391;
   wire N392;
   wire N393;
   wire N394;
   wire N395;
   wire N396;
   wire N397;
   wire N398;
   wire N399;
   wire N400;
   wire N401;
   wire N402;
   wire N403;
   wire N404;
   wire N405;
   wire N406;
   wire N407;
   wire N408;
   wire N409;
   wire N410;
   wire N411;
   wire N412;
   wire N421;
   wire N422;
   wire N423;
   wire N424;
   wire N425;
   wire N426;
   wire N427;
   wire N428;
   wire N429;
   wire N430;
   wire N431;
   wire N432;
   wire N433;
   wire N434;
   wire N435;
   wire N436;
   wire N437;
   wire N438;
   wire N439;
   wire N440;
   wire N441;
   wire N442;
   wire N443;
   wire N444;
   wire n1;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n182;
   wire n368;
   wire n369;
   wire n370;
   wire n371;
   wire n372;
   wire n373;
   wire n374;
   wire n375;
   wire n376;
   wire n377;
   wire n378;
   wire n379;
   wire n380;
   wire n381;
   wire n382;
   wire n383;
   wire n384;
   wire n385;
   wire n386;
   wire n387;
   wire n388;
   wire n389;
   wire n390;
   wire n391;
   wire n392;
   wire n393;
   wire n394;
   wire n395;
   wire n396;
   wire n397;
   wire n398;
   wire n399;
   wire n400;
   wire n401;
   wire n402;
   wire n403;
   wire n404;
   wire n405;
   wire n406;
   wire n407;
   wire n408;
   wire n409;
   wire n410;
   wire n411;
   wire n412;
   wire n413;
   wire n414;
   wire n415;
   wire n416;
   wire n417;
   wire n418;
   wire n419;
   wire n420;
   wire n421;
   wire n422;
   wire n423;
   wire n424;
   wire n425;
   wire n426;
   wire n427;
   wire n428;
   wire n429;
   wire n430;
   wire n431;
   wire n432;
   wire n433;
   wire n434;
   wire n435;
   wire n436;
   wire n437;
   wire n438;
   wire n439;
   wire n440;
   wire n441;
   wire n442;
   wire n443;
   wire n444;
   wire n445;
   wire n446;
   wire n447;
   wire \add_49/carry[5] ;
   wire \add_49/carry[4] ;
   wire \add_49/carry[3] ;
   wire \add_49/carry[2] ;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n179;
   wire n180;
   wire n181;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire [7:0] X6x;
   wire [7:0] X2x;
   wire [7:0] X3x;
   wire [7:0] X7x;
   wire [7:0] X0x;
   wire [7:0] X4x;
   wire [7:0] X5x;
   wire [7:0] X1x;
   wire [7:0] F0X6;
   wire [7:0] F0X2;
   wire [7:0] F0X3;
   wire [7:0] F0X7;
   wire [5:0] i_round;
   wire [7:0] X00x;

   // Module instantiations
   round_funct_DW01_add_0 add_121 (
	.A({ F0X7[7],
		F0X7[6],
		F0X7[5],
		F0X7[4],
		F0X7[3],
		F0X7[2],
		F0X7[1],
		F0X7[0] }),
	.B({ SKx3[7],
		SKx3[6],
		SKx3[5],
		SKx3[4],
		SKx3[3],
		SKx3[2],
		SKx3[1],
		SKx3[0] }),
	.CI(n1),
	.SUM({ N444,
		N443,
		N442,
		N441,
		N440,
		N439,
		N438,
		N437 }));
   round_funct_DW01_sub_0 sub_119 (
	.A({ X6x[7],
		X6x[6],
		X6x[5],
		X6x[4],
		X6x[3],
		X6x[2],
		X6x[1],
		X6x[0] }),
	.B({ N421,
		N422,
		N423,
		N424,
		N425,
		N426,
		N427,
		N428 }),
	.CI(n1),
	.DIFF({ N436,
		N435,
		N434,
		N433,
		N432,
		N431,
		N430,
		N429 }));
   round_funct_DW01_add_1 add_117 (
	.A({ F0X3[7],
		F0X3[6],
		F0X3[5],
		F0X3[4],
		F0X3[3],
		F0X3[2],
		F0X3[1],
		F0X3[0] }),
	.B({ SKx1[7],
		SKx1[6],
		SKx1[5],
		SKx1[4],
		SKx1[3],
		SKx1[2],
		SKx1[1],
		SKx1[0] }),
	.CI(n1),
	.SUM({ N412,
		N411,
		N410,
		N409,
		N408,
		N407,
		N406,
		N405 }));
   round_funct_DW01_sub_1 sub_115 (
	.A({ X2x[7],
		X2x[6],
		X2x[5],
		X2x[4],
		X2x[3],
		X2x[2],
		X2x[1],
		X2x[0] }),
	.B({ N389,
		N390,
		N391,
		N392,
		N393,
		N394,
		N395,
		N396 }),
	.CI(n1),
	.DIFF({ N404,
		N403,
		N402,
		N401,
		N400,
		N399,
		N398,
		N397 }));
   round_funct_DW01_sub_2 sub_106 (
	.A({ X4x[7],
		X4x[6],
		X4x[5],
		X4x[4],
		X4x[3],
		X4x[2],
		X4x[1],
		X4x[0] }),
	.B({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.CI(n1),
	.DIFF({ N302,
		N301,
		N300,
		N299,
		N298,
		N297,
		N296,
		N295 }));
   round_funct_DW01_add_2 add_106 (
	.A({ X4x[7],
		X4x[6],
		X4x[5],
		X4x[4],
		X4x[3],
		X4x[2],
		X4x[1],
		X4x[0] }),
	.B({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.CI(n1),
	.SUM({ N294,
		N293,
		N292,
		N291,
		N290,
		N289,
		N288,
		N287 }));
   round_funct_DW01_sub_3 sub_102 (
	.A({ X0x[7],
		X0x[6],
		X0x[5],
		X0x[4],
		X0x[3],
		X0x[2],
		X0x[1],
		X0x[0] }),
	.B({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.CI(n1),
	.DIFF({ N270,
		N269,
		N268,
		N267,
		N266,
		N265,
		N264,
		N263 }));
   round_funct_DW01_add_3 add_102 (
	.A({ X0x[7],
		X0x[6],
		X0x[5],
		X0x[4],
		X0x[3],
		X0x[2],
		X0x[1],
		X0x[0] }),
	.B({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.CI(n1),
	.SUM({ N262,
		N261,
		N260,
		N259,
		N258,
		N257,
		N256,
		N255 }));
   round_funct_DW01_sub_4 sub_70 (
	.A({ X5x[7],
		X5x[6],
		X5x[5],
		X5x[4],
		X5x[3],
		X5x[2],
		X5x[1],
		X5x[0] }),
	.B({ N14,
		N15,
		N16,
		N17,
		N18,
		N19,
		N20,
		N21 }),
	.CI(n1),
	.DIFF({ N139,
		N138,
		N137,
		N136,
		N135,
		N134,
		N133,
		N132 }));
   round_funct_DW01_sub_5 sub_66 (
	.A({ X1x[7],
		X1x[6],
		X1x[5],
		X1x[4],
		X1x[3],
		X1x[2],
		X1x[1],
		X1x[0] }),
	.B({ N6,
		N7,
		N8,
		N9,
		N10,
		N11,
		N12,
		N13 }),
	.CI(n1),
	.DIFF({ N115,
		N114,
		N113,
		N112,
		N111,
		N110,
		N109,
		N108 }));
   round_funct_DW01_sub_6 sub_57 (
	.A({ P[39],
		P[38],
		P[37],
		P[36],
		P[35],
		P[34],
		P[33],
		P[32] }),
	.B({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.CI(n1),
	.DIFF({ N90,
		N89,
		N88,
		N87,
		N86,
		N85,
		N84,
		N83 }));
   round_funct_DW01_add_4 add_57 (
	.A({ P[39],
		P[38],
		P[37],
		P[36],
		P[35],
		P[34],
		P[33],
		P[32] }),
	.B({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.CI(n1),
	.SUM({ N82,
		N81,
		N80,
		N79,
		N78,
		N77,
		N76,
		N75 }));
   round_funct_DW01_sub_7 sub_53 (
	.A({ P[7],
		P[6],
		P[5],
		P[4],
		P[3],
		P[2],
		P[1],
		P[0] }),
	.B({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.CI(n1),
	.DIFF({ N58,
		N57,
		N56,
		N55,
		N54,
		N53,
		N52,
		N51 }));
   round_funct_DW01_add_5 add_53 (
	.A({ P[7],
		P[6],
		P[5],
		P[4],
		P[3],
		P[2],
		P[1],
		P[0] }),
	.B({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.CI(n1),
	.SUM({ N50,
		N49,
		N48,
		N47,
		N46,
		N45,
		N44,
		N43 }));
   round_funct_DW01_add_6 r138 (
	.A({ X5x[7],
		X5x[6],
		X5x[5],
		X5x[4],
		X5x[3],
		X5x[2],
		X5x[1],
		X5x[0] }),
	.B({ N14,
		N15,
		N16,
		N17,
		N18,
		N19,
		N20,
		N21 }),
	.CI(n1),
	.SUM({ N204,
		N203,
		N202,
		N201,
		N200,
		N199,
		N198,
		N197 }));
   round_funct_DW01_add_7 r137 (
	.A({ X1x[7],
		X1x[6],
		X1x[5],
		X1x[4],
		X1x[3],
		X1x[2],
		X1x[1],
		X1x[0] }),
	.B({ N6,
		N7,
		N8,
		N9,
		N10,
		N11,
		N12,
		N13 }),
	.CI(n1),
	.SUM({ N180,
		N179,
		N178,
		N177,
		N176,
		N175,
		N174,
		N173 }));
   round_funct_DW01_add_8 r136 (
	.A({ F0X6[7],
		F0X6[6],
		F0X6[5],
		F0X6[4],
		F0X6[3],
		F0X6[2],
		F0X6[1],
		F0X6[0] }),
	.B({ SKx3[7],
		SKx3[6],
		SKx3[5],
		SKx3[4],
		SKx3[3],
		SKx3[2],
		SKx3[1],
		SKx3[0] }),
	.CI(n1),
	.SUM({ N147,
		N146,
		N145,
		N144,
		N143,
		N142,
		N141,
		N140 }));
   round_funct_DW01_add_9 r134 (
	.A({ F0X2[7],
		F0X2[6],
		F0X2[5],
		F0X2[4],
		F0X2[3],
		F0X2[2],
		F0X2[1],
		F0X2[0] }),
	.B({ SKx1[7],
		SKx1[6],
		SKx1[5],
		SKx1[4],
		SKx1[3],
		SKx1[2],
		SKx1[1],
		SKx1[0] }),
	.CI(n1),
	.SUM({ N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116 }));
   DFECHD \X00x_reg[7]  (
	.Q(X00x[7]),
	.EB(n315),
	.D(X0x[7]),
	.CK(clk));
   DFECHD \X00x_reg[0]  (
	.Q(X00x[0]),
	.EB(n315),
	.D(X0x[0]),
	.CK(clk));
   DFECHD \X00x_reg[1]  (
	.Q(X00x[1]),
	.EB(n315),
	.D(X0x[1]),
	.CK(clk));
   DFECHD \X00x_reg[2]  (
	.Q(X00x[2]),
	.EB(n315),
	.D(X0x[2]),
	.CK(clk));
   DFECHD \X00x_reg[3]  (
	.Q(X00x[3]),
	.EB(n315),
	.D(X0x[3]),
	.CK(clk));
   DFECHD \X00x_reg[4]  (
	.Q(X00x[4]),
	.EB(n315),
	.D(X0x[4]),
	.CK(clk));
   DFECHD \X00x_reg[5]  (
	.Q(X00x[5]),
	.EB(n315),
	.D(X0x[5]),
	.CK(clk));
   DFECHD \X00x_reg[6]  (
	.Q(X00x[6]),
	.EB(n315),
	.D(X0x[6]),
	.CK(clk));
   QDFFEHD \C0_reg[0]  (
	.Q(C[0]),
	.D(n407),
	.CK(clk));
   QDFFEHD \C0_reg[1]  (
	.Q(C[1]),
	.D(n406),
	.CK(clk));
   QDFFEHD \C0_reg[2]  (
	.Q(C[2]),
	.D(n405),
	.CK(clk));
   QDFFEHD \C0_reg[3]  (
	.Q(C[3]),
	.D(n404),
	.CK(clk));
   QDFFEHD \C0_reg[4]  (
	.Q(C[4]),
	.D(n403),
	.CK(clk));
   QDFFEHD \C0_reg[5]  (
	.Q(C[5]),
	.D(n402),
	.CK(clk));
   QDFFEHD \C0_reg[6]  (
	.Q(C[6]),
	.D(n401),
	.CK(clk));
   QDFFEHD \C0_reg[7]  (
	.Q(C[7]),
	.D(n400),
	.CK(clk));
   QDFFEHD \C4_reg[7]  (
	.Q(C[39]),
	.D(n375),
	.CK(clk));
   QDFFEHD \C4_reg[6]  (
	.Q(C[38]),
	.D(n374),
	.CK(clk));
   QDFFEHD \C4_reg[5]  (
	.Q(C[37]),
	.D(n373),
	.CK(clk));
   QDFFEHD \C4_reg[4]  (
	.Q(C[36]),
	.D(n372),
	.CK(clk));
   QDFFEHD \C4_reg[3]  (
	.Q(C[35]),
	.D(n371),
	.CK(clk));
   QDFFEHD \C4_reg[2]  (
	.Q(C[34]),
	.D(n370),
	.CK(clk));
   QDFFEHD \C4_reg[1]  (
	.Q(C[33]),
	.D(n369),
	.CK(clk));
   QDFFEHD \C4_reg[0]  (
	.Q(C[32]),
	.D(n368),
	.CK(clk));
   DFCLRBEHD \i_round_reg[0]  (
	.RB(n332),
	.QB(n5),
	.Q(n306),
	.LD(N23),
	.D(n5),
	.CK(clk));
   QDFFEHD \X3x_reg[6]  (
	.Q(X3x[6]),
	.D(n377),
	.CK(clk));
   QDFFEHD \X3x_reg[5]  (
	.Q(X3x[5]),
	.D(n378),
	.CK(clk));
   QDFFEHD \X3x_reg[1]  (
	.Q(X3x[1]),
	.D(n382),
	.CK(clk));
   QDFFEHD \X3x_reg[2]  (
	.Q(X3x[2]),
	.D(n381),
	.CK(clk));
   QDFFEHD \X3x_reg[3]  (
	.Q(X3x[3]),
	.D(n380),
	.CK(clk));
   QDFFEHD \X3x_reg[4]  (
	.Q(X3x[4]),
	.D(n379),
	.CK(clk));
   QDFFEHD \X3x_reg[0]  (
	.Q(X3x[0]),
	.D(n383),
	.CK(clk));
   QDFFEHD \X7x_reg[3]  (
	.Q(X7x[3]),
	.D(n420),
	.CK(clk));
   QDFFEHD \X7x_reg[4]  (
	.Q(X7x[4]),
	.D(n419),
	.CK(clk));
   QDFFEHD \X7x_reg[0]  (
	.Q(X7x[0]),
	.D(n423),
	.CK(clk));
   QDFFEHD \X7x_reg[5]  (
	.Q(X7x[5]),
	.D(n418),
	.CK(clk));
   QDFFEHD \X7x_reg[2]  (
	.Q(X7x[2]),
	.D(n421),
	.CK(clk));
   QDFFEHD \X6x_reg[4]  (
	.Q(X6x[4]),
	.D(n427),
	.CK(clk));
   QDFFEHD \X6x_reg[5]  (
	.Q(X6x[5]),
	.D(n426),
	.CK(clk));
   QDFFEHD \X4x_reg[7]  (
	.Q(X4x[7]),
	.D(n439),
	.CK(clk));
   QDFFEHD \X4x_reg[0]  (
	.Q(X4x[0]),
	.D(n446),
	.CK(clk));
   QDFFEHD \X1x_reg[7]  (
	.Q(X1x[7]),
	.D(n392),
	.CK(clk));
   QDFFEHD \X1x_reg[0]  (
	.Q(X1x[0]),
	.D(n399),
	.CK(clk));
   QDFFEHD \X0x_reg[7]  (
	.Q(X0x[7]),
	.D(n408),
	.CK(clk));
   QDFFEHD \X0x_reg[0]  (
	.Q(X0x[0]),
	.D(n415),
	.CK(clk));
   QDFFEHD \X2x_reg[4]  (
	.Q(X2x[4]),
	.D(n387),
	.CK(clk));
   QDFFEHD \X4x_reg[1]  (
	.Q(X4x[1]),
	.D(n445),
	.CK(clk));
   QDFFEHD \X1x_reg[6]  (
	.Q(X1x[6]),
	.D(n393),
	.CK(clk));
   QDFFEHD \X1x_reg[3]  (
	.Q(X1x[3]),
	.D(n396),
	.CK(clk));
   QDFFEHD \X1x_reg[4]  (
	.Q(X1x[4]),
	.D(n395),
	.CK(clk));
   QDFFEHD \X1x_reg[1]  (
	.Q(X1x[1]),
	.D(n398),
	.CK(clk));
   QDFFEHD \X0x_reg[1]  (
	.Q(X0x[1]),
	.D(n414),
	.CK(clk));
   QDFFEHD \X2x_reg[5]  (
	.Q(X2x[5]),
	.D(n386),
	.CK(clk));
   QDFFEHD \X3x_reg[7]  (
	.Q(X3x[7]),
	.D(n376),
	.CK(clk));
   QDFFEHD \X7x_reg[7]  (
	.Q(X7x[7]),
	.D(n416),
	.CK(clk));
   QDFFEHD \X7x_reg[6]  (
	.Q(X7x[6]),
	.D(n417),
	.CK(clk));
   QDFFEHD \X6x_reg[7]  (
	.Q(X6x[7]),
	.D(n424),
	.CK(clk));
   QDFFEHD \X7x_reg[1]  (
	.Q(X7x[1]),
	.D(n422),
	.CK(clk));
   QDFFEHD \X6x_reg[6]  (
	.Q(X6x[6]),
	.D(n425),
	.CK(clk));
   QDFFEHD \X2x_reg[0]  (
	.Q(X2x[0]),
	.D(n391),
	.CK(clk));
   QDFFEHD \X2x_reg[1]  (
	.Q(X2x[1]),
	.D(n390),
	.CK(clk));
   QDFFEHD \X2x_reg[2]  (
	.Q(X2x[2]),
	.D(n389),
	.CK(clk));
   QDFFEHD \X6x_reg[3]  (
	.Q(X6x[3]),
	.D(n428),
	.CK(clk));
   QDFFEHD \X6x_reg[0]  (
	.Q(X6x[0]),
	.D(n431),
	.CK(clk));
   QDFFEHD \X6x_reg[1]  (
	.Q(X6x[1]),
	.D(n430),
	.CK(clk));
   QDFFEHD \X6x_reg[2]  (
	.Q(X6x[2]),
	.D(n429),
	.CK(clk));
   QDFFEHD \X2x_reg[7]  (
	.Q(X2x[7]),
	.D(n384),
	.CK(clk));
   QDFFEHD \X2x_reg[6]  (
	.Q(X2x[6]),
	.D(n385),
	.CK(clk));
   QDFFEHD \X2x_reg[3]  (
	.Q(X2x[3]),
	.D(n388),
	.CK(clk));
   QDFFEHD \X4x_reg[6]  (
	.Q(X4x[6]),
	.D(n440),
	.CK(clk));
   QDFFEHD \X4x_reg[4]  (
	.Q(X4x[4]),
	.D(n442),
	.CK(clk));
   QDFFEHD \X4x_reg[3]  (
	.Q(X4x[3]),
	.D(n443),
	.CK(clk));
   QDFFEHD \X0x_reg[6]  (
	.Q(X0x[6]),
	.D(n409),
	.CK(clk));
   QDFFEHD \X0x_reg[3]  (
	.Q(X0x[3]),
	.D(n412),
	.CK(clk));
   QDFFEHD \X0x_reg[4]  (
	.Q(X0x[4]),
	.D(n411),
	.CK(clk));
   QDFFEHD \X4x_reg[5]  (
	.Q(X4x[5]),
	.D(n441),
	.CK(clk));
   QDFFEHD \X4x_reg[2]  (
	.Q(X4x[2]),
	.D(n444),
	.CK(clk));
   QDFFEHD \X1x_reg[5]  (
	.Q(X1x[5]),
	.D(n394),
	.CK(clk));
   QDFFEHD \X1x_reg[2]  (
	.Q(X1x[2]),
	.D(n397),
	.CK(clk));
   QDFFEHD \X0x_reg[5]  (
	.Q(X0x[5]),
	.D(n410),
	.CK(clk));
   QDFFEHD \X0x_reg[2]  (
	.Q(X0x[2]),
	.D(n413),
	.CK(clk));
   DFECHD \C2_reg[7]  (
	.Q(C[23]),
	.EB(n182),
	.D(n316),
	.CK(clk));
   DFECHD \C6_reg[6]  (
	.Q(C[54]),
	.EB(n182),
	.D(n318),
	.CK(clk));
   DFECHD \C2_reg[0]  (
	.Q(C[16]),
	.EB(n182),
	.D(n319),
	.CK(clk));
   DFECHD \C6_reg[0]  (
	.Q(C[48]),
	.EB(n182),
	.D(n321),
	.CK(clk));
   DFECHD \C6_reg[1]  (
	.Q(C[49]),
	.EB(n182),
	.D(n322),
	.CK(clk));
   DFECHD \C2_reg[1]  (
	.Q(C[17]),
	.EB(n182),
	.D(n323),
	.CK(clk));
   DFECHD \C6_reg[2]  (
	.Q(C[50]),
	.EB(n182),
	.D(n324),
	.CK(clk));
   DFECHD \C2_reg[2]  (
	.Q(C[18]),
	.EB(n182),
	.D(n325),
	.CK(clk));
   DFECHD \C6_reg[3]  (
	.Q(C[51]),
	.EB(n182),
	.D(n326),
	.CK(clk));
   DFECHD \C2_reg[3]  (
	.Q(C[19]),
	.EB(n182),
	.D(n327),
	.CK(clk));
   DFECHD \C6_reg[4]  (
	.Q(C[52]),
	.EB(n182),
	.D(n328),
	.CK(clk));
   DFECHD \C6_reg[7]  (
	.Q(C[55]),
	.EB(n182),
	.D(n329),
	.CK(clk));
   DFECHD \C2_reg[4]  (
	.Q(C[20]),
	.EB(n182),
	.D(n330),
	.CK(clk));
   DFECHD \C2_reg[5]  (
	.Q(C[21]),
	.EB(n182),
	.D(n320),
	.CK(clk));
   DFECHD \C6_reg[5]  (
	.Q(C[53]),
	.EB(n182),
	.D(n331),
	.CK(clk));
   DFECHD \C2_reg[6]  (
	.Q(C[22]),
	.EB(n182),
	.D(n317),
	.CK(clk));
   DFECHD \C3_reg[0]  (
	.Q(C[24]),
	.EB(n182),
	.D(X3x[0]),
	.CK(clk));
   DFECHD \C3_reg[7]  (
	.Q(C[31]),
	.EB(n182),
	.D(X3x[7]),
	.CK(clk));
   DFECHD \C3_reg[6]  (
	.Q(C[30]),
	.EB(n182),
	.D(X3x[6]),
	.CK(clk));
   DFECHD \C7_reg[7]  (
	.Q(C[63]),
	.EB(n182),
	.D(X7x[7]),
	.CK(clk));
   DFECHD \C7_reg[6]  (
	.Q(C[62]),
	.EB(n182),
	.D(X7x[6]),
	.CK(clk));
   DFECHD \C7_reg[0]  (
	.Q(C[56]),
	.EB(n182),
	.D(X7x[0]),
	.CK(clk));
   DFECHD \C1_reg[0]  (
	.Q(C[8]),
	.EB(n182),
	.D(X1x[0]),
	.CK(clk));
   DFECHD \C7_reg[1]  (
	.Q(C[57]),
	.EB(n182),
	.D(X7x[1]),
	.CK(clk));
   DFECHD \C1_reg[1]  (
	.Q(C[9]),
	.EB(n182),
	.D(X1x[1]),
	.CK(clk));
   DFECHD \C3_reg[1]  (
	.Q(C[25]),
	.EB(n182),
	.D(X3x[1]),
	.CK(clk));
   DFECHD \C5_reg[1]  (
	.Q(C[41]),
	.EB(n182),
	.D(X5x[1]),
	.CK(clk));
   DFECHD \C7_reg[2]  (
	.Q(C[58]),
	.EB(n182),
	.D(X7x[2]),
	.CK(clk));
   DFECHD \C1_reg[2]  (
	.Q(C[10]),
	.EB(n182),
	.D(X1x[2]),
	.CK(clk));
   DFECHD \C3_reg[2]  (
	.Q(C[26]),
	.EB(n182),
	.D(X3x[2]),
	.CK(clk));
   DFECHD \C5_reg[2]  (
	.Q(C[42]),
	.EB(n182),
	.D(X5x[2]),
	.CK(clk));
   DFECHD \C7_reg[3]  (
	.Q(C[59]),
	.EB(n182),
	.D(X7x[3]),
	.CK(clk));
   DFECHD \C1_reg[3]  (
	.Q(C[11]),
	.EB(n182),
	.D(X1x[3]),
	.CK(clk));
   DFECHD \C3_reg[3]  (
	.Q(C[27]),
	.EB(n182),
	.D(X3x[3]),
	.CK(clk));
   DFECHD \C5_reg[3]  (
	.Q(C[43]),
	.EB(n182),
	.D(X5x[3]),
	.CK(clk));
   DFECHD \C7_reg[4]  (
	.Q(C[60]),
	.EB(n182),
	.D(X7x[4]),
	.CK(clk));
   DFECHD \C1_reg[4]  (
	.Q(C[12]),
	.EB(n182),
	.D(X1x[4]),
	.CK(clk));
   DFECHD \C3_reg[4]  (
	.Q(C[28]),
	.EB(n182),
	.D(X3x[4]),
	.CK(clk));
   DFECHD \C5_reg[4]  (
	.Q(C[44]),
	.EB(n182),
	.D(X5x[4]),
	.CK(clk));
   DFECHD \C5_reg[5]  (
	.Q(C[45]),
	.EB(n182),
	.D(X5x[5]),
	.CK(clk));
   DFECHD \C3_reg[5]  (
	.Q(C[29]),
	.EB(n182),
	.D(X3x[5]),
	.CK(clk));
   DFECHD \C7_reg[5]  (
	.Q(C[61]),
	.EB(n182),
	.D(X7x[5]),
	.CK(clk));
   DFECHD \C1_reg[5]  (
	.Q(C[13]),
	.EB(n182),
	.D(X1x[5]),
	.CK(clk));
   DFECHD \C1_reg[6]  (
	.Q(C[14]),
	.EB(n182),
	.D(X1x[6]),
	.CK(clk));
   DFECHD \C1_reg[7]  (
	.Q(C[15]),
	.EB(n182),
	.D(X1x[7]),
	.CK(clk));
   DFECHD \C5_reg[6]  (
	.Q(C[46]),
	.EB(n182),
	.D(X5x[6]),
	.CK(clk));
   DFECHD \C5_reg[7]  (
	.Q(C[47]),
	.EB(n182),
	.D(X5x[7]),
	.CK(clk));
   DFECHD \C5_reg[0]  (
	.Q(C[40]),
	.EB(n182),
	.D(X5x[0]),
	.CK(clk));
   DFCLRBEHD \i_round_reg[5]  (
	.RB(n332),
	.QB(n108),
	.Q(i_round[5]),
	.LD(N23),
	.D(N30),
	.CK(clk));
   DFCLRBEHD \i_round_reg[4]  (
	.RB(n332),
	.QB(n104),
	.Q(i_round[4]),
	.LD(N23),
	.D(N29),
	.CK(clk));
   DFCLRBEHD \i_round_reg[3]  (
	.RB(n332),
	.QB(n105),
	.Q(i_round[3]),
	.LD(N23),
	.D(N28),
	.CK(clk));
   DFCLRBEHD \i_round_reg[2]  (
	.RB(n332),
	.QB(n106),
	.Q(i_round[2]),
	.LD(N23),
	.D(N27),
	.CK(clk));
   DFCLRBEHD \i_round_reg[1]  (
	.RB(n332),
	.QB(n107),
	.Q(n311),
	.LD(N23),
	.D(N26),
	.CK(clk));
   DFFCHD \X5x_reg[7]  (
	.QB(n171),
	.Q(X5x[7]),
	.D(n432),
	.CK(clk));
   DFFCHD \X5x_reg[4]  (
	.QB(n174),
	.Q(X5x[4]),
	.D(n435),
	.CK(clk));
   DFFCHD \X5x_reg[3]  (
	.QB(n175),
	.Q(X5x[3]),
	.D(n436),
	.CK(clk));
   DFFCHD \X5x_reg[6]  (
	.QB(n172),
	.Q(X5x[6]),
	.D(n433),
	.CK(clk));
   DFFCHD \X5x_reg[5]  (
	.QB(n173),
	.Q(X5x[5]),
	.D(n434),
	.CK(clk));
   DFFCHD \X5x_reg[1]  (
	.QB(n177),
	.Q(X5x[1]),
	.D(n438),
	.CK(clk));
   DFFCHD \X5x_reg[0]  (
	.QB(n178),
	.Q(X5x[0]),
	.D(n447),
	.CK(clk));
   DFFCHD \X5x_reg[2]  (
	.QB(n176),
	.Q(X5x[2]),
	.D(n437),
	.CK(clk));
   AN3EHD U3 (
	.O(n2),
	.I3(n305),
	.I2(n246),
	.I1(n108));
   OA112EHD U4 (
	.O(n3),
	.C2(n308),
	.C1(n306),
	.B1(n309),
	.A1(n246));
   AN2EHD U5 (
	.O(n4),
	.I2(n309),
	.I1(ed));
   INVDHD U6 (
	.O(n113),
	.I(n162));
   INVDHD U7 (
	.O(n179),
	.I(n112));
   NR2CHD U9 (
	.O(n112),
	.I2(n2),
	.I1(n113));
   NR3BHD U11 (
	.O(n162),
	.I3(n111),
	.I2(n3),
	.I1(n4));
   NR2CHD U44 (
	.O(n247),
	.I2(n182),
	.I1(n246));
   NR2CHD U45 (
	.O(n119),
	.I2(n246),
	.I1(n245));
   NR2CHD U53 (
	.O(n117),
	.I2(ed),
	.I1(n245));
   NR2CHD U55 (
	.O(n248),
	.I2(ed),
	.I1(n182));
   HA1EHD U56 (
	.S(N26),
	.C(\add_49/carry[2] ),
	.B(n306),
	.A(n311));
   HA1EHD U57 (
	.S(N27),
	.C(\add_49/carry[3] ),
	.B(\add_49/carry[2] ),
	.A(i_round[2]));
   HA1EHD U58 (
	.S(N28),
	.C(\add_49/carry[4] ),
	.B(\add_49/carry[3] ),
	.A(i_round[3]));
   HA1EHD U59 (
	.S(N29),
	.C(\add_49/carry[5] ),
	.B(\add_49/carry[4] ),
	.A(i_round[4]));
   TIE0DHD U60 (
	.O(n1));
   XOR2CHD U61 (
	.O(N30),
	.I2(i_round[5]),
	.I1(\add_49/carry[5] ));
   NR2BHD U62 (
	.O(n315),
	.I2(n2),
	.I1(n3));
   XOR2CHD U63 (
	.O(n316),
	.I2(WK1_5[7]),
	.I1(X2x[7]));
   XOR2CHD U64 (
	.O(n317),
	.I2(WK1_5[6]),
	.I1(X2x[6]));
   XOR2CHD U65 (
	.O(n318),
	.I2(WK3_7[6]),
	.I1(X6x[6]));
   XOR2CHD U66 (
	.O(n319),
	.I2(WK1_5[0]),
	.I1(X2x[0]));
   XOR2CHD U67 (
	.O(n320),
	.I2(WK1_5[5]),
	.I1(X2x[5]));
   XOR2CHD U68 (
	.O(n321),
	.I2(WK3_7[0]),
	.I1(X6x[0]));
   XOR2CHD U69 (
	.O(n322),
	.I2(WK3_7[1]),
	.I1(X6x[1]));
   XOR2CHD U70 (
	.O(n323),
	.I2(WK1_5[1]),
	.I1(X2x[1]));
   XOR2CHD U71 (
	.O(n324),
	.I2(WK3_7[2]),
	.I1(X6x[2]));
   XOR2CHD U72 (
	.O(n325),
	.I2(WK1_5[2]),
	.I1(X2x[2]));
   XOR2CHD U73 (
	.O(n326),
	.I2(WK3_7[3]),
	.I1(X6x[3]));
   XOR2CHD U74 (
	.O(n327),
	.I2(WK1_5[3]),
	.I1(X2x[3]));
   XOR2CHD U75 (
	.O(n328),
	.I2(WK3_7[4]),
	.I1(X6x[4]));
   XOR2CHD U76 (
	.O(n329),
	.I2(WK3_7[7]),
	.I1(X6x[7]));
   XOR2CHD U77 (
	.O(n330),
	.I2(WK1_5[4]),
	.I1(X2x[4]));
   XOR2CHD U78 (
	.O(n331),
	.I2(WK3_7[5]),
	.I1(X6x[5]));
   INVCHD U79 (
	.O(n332),
	.I(reset));
   ND2CHD U80 (
	.O(n447),
	.I2(n110),
	.I1(n109));
   AOI222BHD U81 (
	.O(n110),
	.C2(X5x[0]),
	.C1(n112),
	.B2(n2),
	.B1(N132),
	.A2(n111),
	.A1(P[40]));
   AOI22BHD U82 (
	.O(n109),
	.B2(n3),
	.B1(N429),
	.A2(n4),
	.A1(X4x[0]));
   OAI112BHD U83 (
	.O(n446),
	.C2(n114),
	.C1(n113),
	.B1(n116),
	.A1(n115));
   AOI222BHD U84 (
	.O(n116),
	.C2(n119),
	.C1(N75),
	.B2(n118),
	.B1(n4),
	.A2(n117),
	.A1(N83));
   ND2CHD U85 (
	.O(n115),
	.I2(X5x[0]),
	.I1(n3));
   INVCHD U86 (
	.O(n114),
	.I(X4x[0]));
   OAI112BHD U87 (
	.O(n445),
	.C2(n120),
	.C1(n113),
	.B1(n122),
	.A1(n121));
   AOI222BHD U88 (
	.O(n122),
	.C2(n119),
	.C1(N76),
	.B2(n123),
	.B1(n4),
	.A2(n117),
	.A1(N84));
   ND2CHD U89 (
	.O(n121),
	.I2(X5x[1]),
	.I1(n3));
   INVCHD U90 (
	.O(n120),
	.I(X4x[1]));
   OAI112BHD U91 (
	.O(n444),
	.C2(n124),
	.C1(n113),
	.B1(n126),
	.A1(n125));
   AOI222BHD U92 (
	.O(n126),
	.C2(n119),
	.C1(N77),
	.B2(n127),
	.B1(n4),
	.A2(n117),
	.A1(N85));
   ND2CHD U93 (
	.O(n125),
	.I2(X5x[2]),
	.I1(n3));
   INVCHD U94 (
	.O(n124),
	.I(X4x[2]));
   OAI112BHD U95 (
	.O(n443),
	.C2(n128),
	.C1(n113),
	.B1(n130),
	.A1(n129));
   AOI222BHD U96 (
	.O(n130),
	.C2(n119),
	.C1(N78),
	.B2(n131),
	.B1(n4),
	.A2(n117),
	.A1(N86));
   ND2CHD U97 (
	.O(n129),
	.I2(X5x[3]),
	.I1(n3));
   INVCHD U98 (
	.O(n128),
	.I(X4x[3]));
   OAI112BHD U99 (
	.O(n442),
	.C2(n132),
	.C1(n113),
	.B1(n134),
	.A1(n133));
   AOI222BHD U100 (
	.O(n134),
	.C2(n119),
	.C1(N79),
	.B2(n135),
	.B1(n4),
	.A2(n117),
	.A1(N87));
   ND2CHD U101 (
	.O(n133),
	.I2(X5x[4]),
	.I1(n3));
   INVCHD U102 (
	.O(n132),
	.I(X4x[4]));
   OAI112BHD U103 (
	.O(n441),
	.C2(n136),
	.C1(n113),
	.B1(n138),
	.A1(n137));
   AOI222BHD U104 (
	.O(n138),
	.C2(n119),
	.C1(N80),
	.B2(n139),
	.B1(n4),
	.A2(n117),
	.A1(N88));
   ND2CHD U105 (
	.O(n137),
	.I2(X5x[5]),
	.I1(n3));
   INVCHD U106 (
	.O(n136),
	.I(X4x[5]));
   OAI112BHD U107 (
	.O(n440),
	.C2(n140),
	.C1(n113),
	.B1(n142),
	.A1(n141));
   AOI222BHD U108 (
	.O(n142),
	.C2(n119),
	.C1(N81),
	.B2(n143),
	.B1(n4),
	.A2(n117),
	.A1(N89));
   ND2CHD U109 (
	.O(n141),
	.I2(X5x[6]),
	.I1(n3));
   INVCHD U110 (
	.O(n140),
	.I(X4x[6]));
   OAI112BHD U111 (
	.O(n439),
	.C2(n144),
	.C1(n113),
	.B1(n146),
	.A1(n145));
   AOI222BHD U112 (
	.O(n146),
	.C2(n119),
	.C1(N82),
	.B2(n147),
	.B1(n4),
	.A2(n117),
	.A1(N90));
   ND2CHD U113 (
	.O(n145),
	.I2(X5x[7]),
	.I1(n3));
   INVCHD U114 (
	.O(n144),
	.I(X4x[7]));
   ND2CHD U115 (
	.O(n438),
	.I2(n149),
	.I1(n148));
   AOI222BHD U116 (
	.O(n149),
	.C2(X5x[1]),
	.C1(n112),
	.B2(n2),
	.B1(N133),
	.A2(n111),
	.A1(P[41]));
   AOI22BHD U117 (
	.O(n148),
	.B2(n3),
	.B1(N430),
	.A2(n4),
	.A1(X4x[1]));
   ND2CHD U118 (
	.O(n437),
	.I2(n151),
	.I1(n150));
   AOI222BHD U119 (
	.O(n151),
	.C2(X5x[2]),
	.C1(n112),
	.B2(n2),
	.B1(N134),
	.A2(n111),
	.A1(P[42]));
   AOI22BHD U120 (
	.O(n150),
	.B2(n3),
	.B1(N431),
	.A2(n4),
	.A1(X4x[2]));
   ND2CHD U121 (
	.O(n436),
	.I2(n153),
	.I1(n152));
   AOI222BHD U122 (
	.O(n153),
	.C2(X5x[3]),
	.C1(n112),
	.B2(n2),
	.B1(N135),
	.A2(n111),
	.A1(P[43]));
   AOI22BHD U123 (
	.O(n152),
	.B2(n3),
	.B1(N432),
	.A2(n4),
	.A1(X4x[3]));
   ND2CHD U124 (
	.O(n435),
	.I2(n155),
	.I1(n154));
   AOI222BHD U125 (
	.O(n155),
	.C2(X5x[4]),
	.C1(n112),
	.B2(n2),
	.B1(N136),
	.A2(n111),
	.A1(P[44]));
   AOI22BHD U126 (
	.O(n154),
	.B2(n3),
	.B1(N433),
	.A2(n4),
	.A1(X4x[4]));
   ND2CHD U127 (
	.O(n434),
	.I2(n157),
	.I1(n156));
   AOI222BHD U128 (
	.O(n157),
	.C2(X5x[5]),
	.C1(n112),
	.B2(n2),
	.B1(N137),
	.A2(n111),
	.A1(P[45]));
   AOI22BHD U129 (
	.O(n156),
	.B2(n3),
	.B1(N434),
	.A2(n4),
	.A1(X4x[5]));
   ND2CHD U130 (
	.O(n433),
	.I2(n159),
	.I1(n158));
   AOI222BHD U131 (
	.O(n159),
	.C2(X5x[6]),
	.C1(n112),
	.B2(n2),
	.B1(N138),
	.A2(n111),
	.A1(P[46]));
   AOI22BHD U132 (
	.O(n158),
	.B2(n3),
	.B1(N435),
	.A2(n4),
	.A1(X4x[6]));
   ND2CHD U133 (
	.O(n432),
	.I2(n161),
	.I1(n160));
   AOI222BHD U134 (
	.O(n161),
	.C2(X5x[7]),
	.C1(n112),
	.B2(n2),
	.B1(N139),
	.A2(n111),
	.A1(P[47]));
   AOI22BHD U135 (
	.O(n160),
	.B2(n3),
	.B1(N436),
	.A2(n4),
	.A1(X4x[7]));
   AO2222BHD U136 (
	.O(n431),
	.D2(n163),
	.D1(n111),
	.C2(X6x[0]),
	.C1(n162),
	.B2(n4),
	.B1(N197),
	.A2(n3),
	.A1(X7x[0]));
   XOR2CHD U137 (
	.O(n163),
	.I2(P[48]),
	.I1(WK3_7[0]));
   AO2222BHD U138 (
	.O(n430),
	.D2(n164),
	.D1(n111),
	.C2(X6x[1]),
	.C1(n162),
	.B2(n4),
	.B1(N198),
	.A2(n3),
	.A1(X7x[1]));
   XOR2CHD U139 (
	.O(n164),
	.I2(P[49]),
	.I1(WK3_7[1]));
   AO2222BHD U140 (
	.O(n429),
	.D2(n165),
	.D1(n111),
	.C2(X6x[2]),
	.C1(n162),
	.B2(n4),
	.B1(N199),
	.A2(n3),
	.A1(X7x[2]));
   XOR2CHD U141 (
	.O(n165),
	.I2(P[50]),
	.I1(WK3_7[2]));
   AO2222BHD U142 (
	.O(n428),
	.D2(n166),
	.D1(n111),
	.C2(X6x[3]),
	.C1(n162),
	.B2(n4),
	.B1(N200),
	.A2(n3),
	.A1(X7x[3]));
   XOR2CHD U143 (
	.O(n166),
	.I2(P[51]),
	.I1(WK3_7[3]));
   AO2222BHD U144 (
	.O(n427),
	.D2(n167),
	.D1(n111),
	.C2(X6x[4]),
	.C1(n162),
	.B2(n4),
	.B1(N201),
	.A2(n3),
	.A1(X7x[4]));
   XOR2CHD U145 (
	.O(n167),
	.I2(P[52]),
	.I1(WK3_7[4]));
   AO2222BHD U146 (
	.O(n426),
	.D2(n168),
	.D1(n111),
	.C2(X6x[5]),
	.C1(n162),
	.B2(n4),
	.B1(N202),
	.A2(n3),
	.A1(X7x[5]));
   XOR2CHD U147 (
	.O(n168),
	.I2(P[53]),
	.I1(WK3_7[5]));
   AO2222BHD U148 (
	.O(n425),
	.D2(n169),
	.D1(n111),
	.C2(X6x[6]),
	.C1(n162),
	.B2(n4),
	.B1(N203),
	.A2(n3),
	.A1(X7x[6]));
   XOR2CHD U149 (
	.O(n169),
	.I2(P[54]),
	.I1(WK3_7[6]));
   AO2222BHD U150 (
	.O(n424),
	.D2(n170),
	.D1(n111),
	.C2(X6x[7]),
	.C1(n162),
	.B2(n4),
	.B1(N204),
	.A2(n3),
	.A1(X7x[7]));
   XOR2CHD U151 (
	.O(n170),
	.I2(P[55]),
	.I1(WK3_7[7]));
   OAI112BHD U152 (
	.O(n423),
	.C2(n180),
	.C1(n179),
	.B1(n183),
	.A1(n181));
   AOI22BHD U153 (
	.O(n183),
	.B2(X6x[0]),
	.B1(n4),
	.A2(n111),
	.A1(P[56]));
   AOI22BHD U154 (
	.O(n181),
	.B2(n2),
	.B1(n185),
	.A2(n3),
	.A1(n184));
   XOR2CHD U155 (
	.O(n184),
	.I2(N437),
	.I1(X00x[0]));
   INVCHD U156 (
	.O(n180),
	.I(X7x[0]));
   OAI112BHD U157 (
	.O(n422),
	.C2(n186),
	.C1(n179),
	.B1(n188),
	.A1(n187));
   AOI22BHD U158 (
	.O(n188),
	.B2(X6x[1]),
	.B1(n4),
	.A2(n111),
	.A1(P[57]));
   AOI22BHD U159 (
	.O(n187),
	.B2(n2),
	.B1(n190),
	.A2(n3),
	.A1(n189));
   XOR2CHD U160 (
	.O(n189),
	.I2(N438),
	.I1(X00x[1]));
   INVCHD U161 (
	.O(n186),
	.I(X7x[1]));
   OAI112BHD U162 (
	.O(n421),
	.C2(n191),
	.C1(n179),
	.B1(n193),
	.A1(n192));
   AOI22BHD U163 (
	.O(n193),
	.B2(X6x[2]),
	.B1(n4),
	.A2(n111),
	.A1(P[58]));
   AOI22BHD U164 (
	.O(n192),
	.B2(n2),
	.B1(n195),
	.A2(n3),
	.A1(n194));
   XOR2CHD U165 (
	.O(n194),
	.I2(N439),
	.I1(X00x[2]));
   INVCHD U166 (
	.O(n191),
	.I(X7x[2]));
   OAI112BHD U167 (
	.O(n420),
	.C2(n196),
	.C1(n179),
	.B1(n198),
	.A1(n197));
   AOI22BHD U168 (
	.O(n198),
	.B2(X6x[3]),
	.B1(n4),
	.A2(n111),
	.A1(P[59]));
   AOI22BHD U169 (
	.O(n197),
	.B2(n2),
	.B1(n200),
	.A2(n3),
	.A1(n199));
   XOR2CHD U170 (
	.O(n199),
	.I2(N440),
	.I1(X00x[3]));
   INVCHD U171 (
	.O(n196),
	.I(X7x[3]));
   OAI112BHD U172 (
	.O(n419),
	.C2(n201),
	.C1(n179),
	.B1(n203),
	.A1(n202));
   AOI22BHD U173 (
	.O(n203),
	.B2(X6x[4]),
	.B1(n4),
	.A2(n111),
	.A1(P[60]));
   AOI22BHD U174 (
	.O(n202),
	.B2(n2),
	.B1(n205),
	.A2(n3),
	.A1(n204));
   XOR2CHD U175 (
	.O(n204),
	.I2(N441),
	.I1(X00x[4]));
   INVCHD U176 (
	.O(n201),
	.I(X7x[4]));
   OAI112BHD U177 (
	.O(n418),
	.C2(n206),
	.C1(n179),
	.B1(n208),
	.A1(n207));
   AOI22BHD U178 (
	.O(n208),
	.B2(X6x[5]),
	.B1(n4),
	.A2(n111),
	.A1(P[61]));
   AOI22BHD U179 (
	.O(n207),
	.B2(n2),
	.B1(n210),
	.A2(n3),
	.A1(n209));
   XOR2CHD U180 (
	.O(n209),
	.I2(N442),
	.I1(X00x[5]));
   INVCHD U181 (
	.O(n206),
	.I(X7x[5]));
   OAI112BHD U182 (
	.O(n417),
	.C2(n211),
	.C1(n179),
	.B1(n213),
	.A1(n212));
   AOI22BHD U183 (
	.O(n213),
	.B2(X6x[6]),
	.B1(n4),
	.A2(n111),
	.A1(P[62]));
   AOI22BHD U184 (
	.O(n212),
	.B2(n2),
	.B1(n215),
	.A2(n3),
	.A1(n214));
   XOR2CHD U185 (
	.O(n214),
	.I2(N443),
	.I1(X00x[6]));
   INVCHD U186 (
	.O(n211),
	.I(X7x[6]));
   OAI112BHD U187 (
	.O(n416),
	.C2(n216),
	.C1(n179),
	.B1(n218),
	.A1(n217));
   AOI22BHD U188 (
	.O(n218),
	.B2(X6x[7]),
	.B1(n4),
	.A2(n111),
	.A1(P[63]));
   AOI22BHD U189 (
	.O(n217),
	.B2(n2),
	.B1(n220),
	.A2(n3),
	.A1(n219));
   XOR2CHD U190 (
	.O(n219),
	.I2(N444),
	.I1(X00x[7]));
   INVCHD U191 (
	.O(n216),
	.I(X7x[7]));
   OAI112BHD U192 (
	.O(n415),
	.C2(n221),
	.C1(n113),
	.B1(n223),
	.A1(n222));
   AOI222BHD U193 (
	.O(n223),
	.C2(n119),
	.C1(N43),
	.B2(n185),
	.B1(n4),
	.A2(n117),
	.A1(N51));
   XOR2CHD U194 (
	.O(n185),
	.I2(N140),
	.I1(X7x[0]));
   ND2CHD U195 (
	.O(n222),
	.I2(n3),
	.I1(X1x[0]));
   INVCHD U196 (
	.O(n221),
	.I(X0x[0]));
   OAI112BHD U197 (
	.O(n414),
	.C2(n224),
	.C1(n113),
	.B1(n226),
	.A1(n225));
   AOI222BHD U198 (
	.O(n226),
	.C2(n119),
	.C1(N44),
	.B2(n190),
	.B1(n4),
	.A2(n117),
	.A1(N52));
   XOR2CHD U199 (
	.O(n190),
	.I2(N141),
	.I1(X7x[1]));
   ND2CHD U200 (
	.O(n225),
	.I2(n3),
	.I1(X1x[1]));
   INVCHD U201 (
	.O(n224),
	.I(X0x[1]));
   OAI112BHD U202 (
	.O(n413),
	.C2(n227),
	.C1(n113),
	.B1(n229),
	.A1(n228));
   AOI222BHD U203 (
	.O(n229),
	.C2(n119),
	.C1(N45),
	.B2(n195),
	.B1(n4),
	.A2(n117),
	.A1(N53));
   XOR2CHD U204 (
	.O(n195),
	.I2(N142),
	.I1(X7x[2]));
   ND2CHD U205 (
	.O(n228),
	.I2(n3),
	.I1(X1x[2]));
   INVCHD U206 (
	.O(n227),
	.I(X0x[2]));
   OAI112BHD U207 (
	.O(n412),
	.C2(n230),
	.C1(n113),
	.B1(n232),
	.A1(n231));
   AOI222BHD U208 (
	.O(n232),
	.C2(n119),
	.C1(N46),
	.B2(n200),
	.B1(n4),
	.A2(n117),
	.A1(N54));
   XOR2CHD U209 (
	.O(n200),
	.I2(N143),
	.I1(X7x[3]));
   ND2CHD U210 (
	.O(n231),
	.I2(n3),
	.I1(X1x[3]));
   INVCHD U211 (
	.O(n230),
	.I(X0x[3]));
   OAI112BHD U212 (
	.O(n411),
	.C2(n233),
	.C1(n113),
	.B1(n235),
	.A1(n234));
   AOI222BHD U213 (
	.O(n235),
	.C2(n119),
	.C1(N47),
	.B2(n205),
	.B1(n4),
	.A2(n117),
	.A1(N55));
   XOR2CHD U214 (
	.O(n205),
	.I2(N144),
	.I1(X7x[4]));
   ND2CHD U215 (
	.O(n234),
	.I2(n3),
	.I1(X1x[4]));
   INVCHD U216 (
	.O(n233),
	.I(X0x[4]));
   OAI112BHD U217 (
	.O(n410),
	.C2(n236),
	.C1(n113),
	.B1(n238),
	.A1(n237));
   AOI222BHD U218 (
	.O(n238),
	.C2(n119),
	.C1(N48),
	.B2(n210),
	.B1(n4),
	.A2(n117),
	.A1(N56));
   XOR2CHD U219 (
	.O(n210),
	.I2(N145),
	.I1(X7x[5]));
   ND2CHD U220 (
	.O(n237),
	.I2(n3),
	.I1(X1x[5]));
   INVCHD U221 (
	.O(n236),
	.I(X0x[5]));
   OAI112BHD U222 (
	.O(n409),
	.C2(n239),
	.C1(n113),
	.B1(n241),
	.A1(n240));
   AOI222BHD U223 (
	.O(n241),
	.C2(n119),
	.C1(N49),
	.B2(n215),
	.B1(n4),
	.A2(n117),
	.A1(N57));
   XOR2CHD U224 (
	.O(n215),
	.I2(N146),
	.I1(X7x[6]));
   ND2CHD U225 (
	.O(n240),
	.I2(n3),
	.I1(X1x[6]));
   INVCHD U226 (
	.O(n239),
	.I(X0x[6]));
   OAI112BHD U227 (
	.O(n408),
	.C2(n242),
	.C1(n113),
	.B1(n244),
	.A1(n243));
   AOI222BHD U228 (
	.O(n244),
	.C2(n119),
	.C1(N50),
	.B2(n220),
	.B1(n4),
	.A2(n117),
	.A1(N58));
   XOR2CHD U229 (
	.O(n220),
	.I2(N147),
	.I1(X7x[7]));
   ND2CHD U230 (
	.O(n243),
	.I2(n3),
	.I1(X1x[7]));
   INVCHD U231 (
	.O(n242),
	.I(X0x[7]));
   AO222CHD U232 (
	.O(n407),
	.C2(n182),
	.C1(C[0]),
	.B2(n248),
	.B1(N263),
	.A2(n247),
	.A1(N255));
   AO222CHD U233 (
	.O(n406),
	.C2(n182),
	.C1(C[1]),
	.B2(n248),
	.B1(N264),
	.A2(n247),
	.A1(N256));
   AO222CHD U234 (
	.O(n405),
	.C2(n182),
	.C1(C[2]),
	.B2(n248),
	.B1(N265),
	.A2(n247),
	.A1(N257));
   AO222CHD U235 (
	.O(n404),
	.C2(n182),
	.C1(C[3]),
	.B2(n248),
	.B1(N266),
	.A2(n247),
	.A1(N258));
   AO222CHD U236 (
	.O(n403),
	.C2(n182),
	.C1(C[4]),
	.B2(n248),
	.B1(N267),
	.A2(n247),
	.A1(N259));
   AO222CHD U237 (
	.O(n402),
	.C2(n182),
	.C1(C[5]),
	.B2(n248),
	.B1(N268),
	.A2(n247),
	.A1(N260));
   AO222CHD U238 (
	.O(n401),
	.C2(n182),
	.C1(C[6]),
	.B2(n248),
	.B1(N269),
	.A2(n247),
	.A1(N261));
   AO222CHD U239 (
	.O(n400),
	.C2(n182),
	.C1(C[7]),
	.B2(n248),
	.B1(N270),
	.A2(n247),
	.A1(N262));
   ND2CHD U240 (
	.O(n399),
	.I2(n250),
	.I1(n249));
   AOI222BHD U241 (
	.O(n250),
	.C2(n112),
	.C1(X1x[0]),
	.B2(n2),
	.B1(N108),
	.A2(n111),
	.A1(P[8]));
   AOI22BHD U242 (
	.O(n249),
	.B2(n3),
	.B1(N397),
	.A2(n4),
	.A1(X0x[0]));
   ND2CHD U243 (
	.O(n398),
	.I2(n252),
	.I1(n251));
   AOI222BHD U244 (
	.O(n252),
	.C2(n112),
	.C1(X1x[1]),
	.B2(n2),
	.B1(N109),
	.A2(n111),
	.A1(P[9]));
   AOI22BHD U245 (
	.O(n251),
	.B2(n3),
	.B1(N398),
	.A2(n4),
	.A1(X0x[1]));
   ND2CHD U246 (
	.O(n397),
	.I2(n254),
	.I1(n253));
   AOI222BHD U247 (
	.O(n254),
	.C2(n112),
	.C1(X1x[2]),
	.B2(n2),
	.B1(N110),
	.A2(n111),
	.A1(P[10]));
   AOI22BHD U248 (
	.O(n253),
	.B2(n3),
	.B1(N399),
	.A2(n4),
	.A1(X0x[2]));
   ND2CHD U249 (
	.O(n396),
	.I2(n256),
	.I1(n255));
   AOI222BHD U250 (
	.O(n256),
	.C2(n112),
	.C1(X1x[3]),
	.B2(n2),
	.B1(N111),
	.A2(n111),
	.A1(P[11]));
   AOI22BHD U251 (
	.O(n255),
	.B2(n3),
	.B1(N400),
	.A2(n4),
	.A1(X0x[3]));
   ND2CHD U252 (
	.O(n395),
	.I2(n258),
	.I1(n257));
   AOI222BHD U253 (
	.O(n258),
	.C2(n112),
	.C1(X1x[4]),
	.B2(n2),
	.B1(N112),
	.A2(n111),
	.A1(P[12]));
   AOI22BHD U254 (
	.O(n257),
	.B2(n3),
	.B1(N401),
	.A2(n4),
	.A1(X0x[4]));
   ND2CHD U255 (
	.O(n394),
	.I2(n260),
	.I1(n259));
   AOI222BHD U256 (
	.O(n260),
	.C2(n112),
	.C1(X1x[5]),
	.B2(n2),
	.B1(N113),
	.A2(n111),
	.A1(P[13]));
   AOI22BHD U257 (
	.O(n259),
	.B2(n3),
	.B1(N402),
	.A2(n4),
	.A1(X0x[5]));
   ND2CHD U258 (
	.O(n393),
	.I2(n262),
	.I1(n261));
   AOI222BHD U259 (
	.O(n262),
	.C2(n112),
	.C1(X1x[6]),
	.B2(n2),
	.B1(N114),
	.A2(n111),
	.A1(P[14]));
   AOI22BHD U260 (
	.O(n261),
	.B2(n3),
	.B1(N403),
	.A2(n4),
	.A1(X0x[6]));
   ND2CHD U261 (
	.O(n392),
	.I2(n264),
	.I1(n263));
   AOI222BHD U262 (
	.O(n264),
	.C2(n112),
	.C1(X1x[7]),
	.B2(n2),
	.B1(N115),
	.A2(n111),
	.A1(P[15]));
   AOI22BHD U263 (
	.O(n263),
	.B2(n3),
	.B1(N404),
	.A2(n4),
	.A1(X0x[7]));
   AO2222BHD U264 (
	.O(n391),
	.D2(n265),
	.D1(n111),
	.C2(X2x[0]),
	.C1(n162),
	.B2(n4),
	.B1(N173),
	.A2(n3),
	.A1(X3x[0]));
   XOR2CHD U265 (
	.O(n265),
	.I2(P[16]),
	.I1(WK1_5[0]));
   AO2222BHD U266 (
	.O(n390),
	.D2(n266),
	.D1(n111),
	.C2(X2x[1]),
	.C1(n162),
	.B2(n4),
	.B1(N174),
	.A2(n3),
	.A1(X3x[1]));
   XOR2CHD U267 (
	.O(n266),
	.I2(P[17]),
	.I1(WK1_5[1]));
   AO2222BHD U268 (
	.O(n389),
	.D2(n267),
	.D1(n111),
	.C2(X2x[2]),
	.C1(n162),
	.B2(n4),
	.B1(N175),
	.A2(n3),
	.A1(X3x[2]));
   XOR2CHD U269 (
	.O(n267),
	.I2(P[18]),
	.I1(WK1_5[2]));
   AO2222BHD U270 (
	.O(n388),
	.D2(n268),
	.D1(n111),
	.C2(X2x[3]),
	.C1(n162),
	.B2(n4),
	.B1(N176),
	.A2(n3),
	.A1(X3x[3]));
   XOR2CHD U271 (
	.O(n268),
	.I2(P[19]),
	.I1(WK1_5[3]));
   AO2222BHD U272 (
	.O(n387),
	.D2(n269),
	.D1(n111),
	.C2(X2x[4]),
	.C1(n162),
	.B2(n4),
	.B1(N177),
	.A2(n3),
	.A1(X3x[4]));
   XOR2CHD U273 (
	.O(n269),
	.I2(P[20]),
	.I1(WK1_5[4]));
   AO2222BHD U274 (
	.O(n386),
	.D2(n270),
	.D1(n111),
	.C2(X2x[5]),
	.C1(n162),
	.B2(n4),
	.B1(N178),
	.A2(n3),
	.A1(X3x[5]));
   XOR2CHD U275 (
	.O(n270),
	.I2(P[21]),
	.I1(WK1_5[5]));
   AO2222BHD U276 (
	.O(n385),
	.D2(n271),
	.D1(n111),
	.C2(X2x[6]),
	.C1(n162),
	.B2(n4),
	.B1(N179),
	.A2(n3),
	.A1(X3x[6]));
   XOR2CHD U277 (
	.O(n271),
	.I2(P[22]),
	.I1(WK1_5[6]));
   AO2222BHD U278 (
	.O(n384),
	.D2(n272),
	.D1(n111),
	.C2(X2x[7]),
	.C1(n162),
	.B2(n4),
	.B1(N180),
	.A2(n3),
	.A1(X3x[7]));
   XOR2CHD U279 (
	.O(n272),
	.I2(P[23]),
	.I1(WK1_5[7]));
   OAI112BHD U280 (
	.O(n383),
	.C2(n273),
	.C1(n179),
	.B1(n275),
	.A1(n274));
   AOI22BHD U281 (
	.O(n275),
	.B2(X2x[0]),
	.B1(n4),
	.A2(n111),
	.A1(P[24]));
   AOI22BHD U282 (
	.O(n274),
	.B2(n2),
	.B1(n118),
	.A2(n276),
	.A1(n3));
   XOR2CHD U283 (
	.O(n118),
	.I2(N116),
	.I1(X3x[0]));
   XOR2CHD U284 (
	.O(n276),
	.I2(N405),
	.I1(X4x[0]));
   INVCHD U285 (
	.O(n273),
	.I(X3x[0]));
   OAI112BHD U286 (
	.O(n382),
	.C2(n277),
	.C1(n179),
	.B1(n279),
	.A1(n278));
   AOI22BHD U287 (
	.O(n279),
	.B2(X2x[1]),
	.B1(n4),
	.A2(n111),
	.A1(P[25]));
   AOI22BHD U288 (
	.O(n278),
	.B2(n2),
	.B1(n123),
	.A2(n280),
	.A1(n3));
   XOR2CHD U289 (
	.O(n123),
	.I2(N117),
	.I1(X3x[1]));
   XOR2CHD U290 (
	.O(n280),
	.I2(N406),
	.I1(X4x[1]));
   INVCHD U291 (
	.O(n277),
	.I(X3x[1]));
   OAI112BHD U292 (
	.O(n381),
	.C2(n281),
	.C1(n179),
	.B1(n283),
	.A1(n282));
   AOI22BHD U293 (
	.O(n283),
	.B2(X2x[2]),
	.B1(n4),
	.A2(n111),
	.A1(P[26]));
   AOI22BHD U294 (
	.O(n282),
	.B2(n2),
	.B1(n127),
	.A2(n284),
	.A1(n3));
   XOR2CHD U295 (
	.O(n127),
	.I2(N118),
	.I1(X3x[2]));
   XOR2CHD U296 (
	.O(n284),
	.I2(N407),
	.I1(X4x[2]));
   INVCHD U297 (
	.O(n281),
	.I(X3x[2]));
   OAI112BHD U298 (
	.O(n380),
	.C2(n285),
	.C1(n179),
	.B1(n287),
	.A1(n286));
   AOI22BHD U299 (
	.O(n287),
	.B2(X2x[3]),
	.B1(n4),
	.A2(n111),
	.A1(P[27]));
   AOI22BHD U300 (
	.O(n286),
	.B2(n2),
	.B1(n131),
	.A2(n288),
	.A1(n3));
   XOR2CHD U301 (
	.O(n131),
	.I2(N119),
	.I1(X3x[3]));
   XOR2CHD U302 (
	.O(n288),
	.I2(N408),
	.I1(X4x[3]));
   INVCHD U303 (
	.O(n285),
	.I(X3x[3]));
   OAI112BHD U304 (
	.O(n379),
	.C2(n289),
	.C1(n179),
	.B1(n291),
	.A1(n290));
   AOI22BHD U305 (
	.O(n291),
	.B2(X2x[4]),
	.B1(n4),
	.A2(n111),
	.A1(P[28]));
   AOI22BHD U306 (
	.O(n290),
	.B2(n2),
	.B1(n135),
	.A2(n292),
	.A1(n3));
   XOR2CHD U307 (
	.O(n135),
	.I2(N120),
	.I1(X3x[4]));
   XOR2CHD U308 (
	.O(n292),
	.I2(N409),
	.I1(X4x[4]));
   INVCHD U309 (
	.O(n289),
	.I(X3x[4]));
   OAI112BHD U310 (
	.O(n378),
	.C2(n293),
	.C1(n179),
	.B1(n295),
	.A1(n294));
   AOI22BHD U311 (
	.O(n295),
	.B2(X2x[5]),
	.B1(n4),
	.A2(n111),
	.A1(P[29]));
   AOI22BHD U312 (
	.O(n294),
	.B2(n2),
	.B1(n139),
	.A2(n296),
	.A1(n3));
   XOR2CHD U313 (
	.O(n139),
	.I2(N121),
	.I1(X3x[5]));
   XOR2CHD U314 (
	.O(n296),
	.I2(N410),
	.I1(X4x[5]));
   INVCHD U315 (
	.O(n293),
	.I(X3x[5]));
   OAI112BHD U316 (
	.O(n377),
	.C2(n297),
	.C1(n179),
	.B1(n299),
	.A1(n298));
   AOI22BHD U317 (
	.O(n299),
	.B2(X2x[6]),
	.B1(n4),
	.A2(n111),
	.A1(P[30]));
   AOI22BHD U318 (
	.O(n298),
	.B2(n2),
	.B1(n143),
	.A2(n300),
	.A1(n3));
   XOR2CHD U319 (
	.O(n143),
	.I2(N122),
	.I1(X3x[6]));
   XOR2CHD U320 (
	.O(n300),
	.I2(N411),
	.I1(X4x[6]));
   INVCHD U321 (
	.O(n297),
	.I(X3x[6]));
   OAI112BHD U322 (
	.O(n376),
	.C2(n301),
	.C1(n179),
	.B1(n303),
	.A1(n302));
   AOI22BHD U323 (
	.O(n303),
	.B2(X2x[7]),
	.B1(n4),
	.A2(n111),
	.A1(P[31]));
   AOI22BHD U324 (
	.O(n302),
	.B2(n2),
	.B1(n147),
	.A2(n304),
	.A1(n3));
   XOR2CHD U325 (
	.O(n147),
	.I2(N123),
	.I1(X3x[7]));
   XOR2CHD U326 (
	.O(n304),
	.I2(N412),
	.I1(X4x[7]));
   INVCHD U327 (
	.O(n301),
	.I(X3x[7]));
   INVDHD U328 (
	.O(n111),
	.I(n245));
   ND3CHD U329 (
	.O(n245),
	.I3(n307),
	.I2(n306),
	.I1(n108));
   OR2B1CHD U330 (
	.O(n308),
	.I1(n310),
	.B1(n108));
   XOR2CHD U331 (
	.O(n309),
	.I2(n307),
	.I1(n108));
   NR2BHD U332 (
	.O(n307),
	.I2(n310),
	.I1(n311));
   AO222CHD U333 (
	.O(n375),
	.C2(n182),
	.C1(C[39]),
	.B2(n248),
	.B1(N302),
	.A2(n247),
	.A1(N294));
   AO222CHD U334 (
	.O(n374),
	.C2(n182),
	.C1(C[38]),
	.B2(n248),
	.B1(N301),
	.A2(n247),
	.A1(N293));
   AO222CHD U335 (
	.O(n373),
	.C2(n182),
	.C1(C[37]),
	.B2(n248),
	.B1(N300),
	.A2(n247),
	.A1(N292));
   AO222CHD U336 (
	.O(n372),
	.C2(n182),
	.C1(C[36]),
	.B2(n248),
	.B1(N299),
	.A2(n247),
	.A1(N291));
   AO222CHD U337 (
	.O(n371),
	.C2(n182),
	.C1(C[35]),
	.B2(n248),
	.B1(N298),
	.A2(n247),
	.A1(N290));
   AO222CHD U338 (
	.O(n370),
	.C2(n182),
	.C1(C[34]),
	.B2(n248),
	.B1(N297),
	.A2(n247),
	.A1(N289));
   AO222CHD U339 (
	.O(n369),
	.C2(n182),
	.C1(C[33]),
	.B2(n248),
	.B1(N296),
	.A2(n247),
	.A1(N288));
   AO222CHD U340 (
	.O(n368),
	.C2(n182),
	.C1(C[32]),
	.B2(n248),
	.B1(N295),
	.A2(n247),
	.A1(N287));
   INVCHD U341 (
	.O(n246),
	.I(ed));
   ND2HHD U342 (
	.O(n182),
	.I2(i_round[5]),
	.I1(n305));
   NR3BHD U343 (
	.O(n305),
	.I3(n306),
	.I2(n107),
	.I1(n310));
   XOR4EHD U344 (
	.O(N9),
	.I4(X0x[1]),
	.I3(X0x[6]),
	.I2(SKx0[4]),
	.I1(X0x[0]));
   XOR4EHD U345 (
	.O(N8),
	.I4(X0x[2]),
	.I3(X0x[7]),
	.I2(SKx0[5]),
	.I1(X0x[1]));
   XOR4EHD U346 (
	.O(N7),
	.I4(X0x[2]),
	.I3(X0x[3]),
	.I2(SKx0[6]),
	.I1(X0x[0]));
   XOR4EHD U347 (
	.O(N6),
	.I4(X0x[3]),
	.I3(X0x[4]),
	.I2(SKx0[7]),
	.I1(X0x[1]));
   XOR4EHD U348 (
	.O(N428),
	.I4(n173),
	.I3(SKx2[0]),
	.I2(X5x[4]),
	.I1(n176));
   XOR4EHD U349 (
	.O(N427),
	.I4(n172),
	.I3(SKx2[1]),
	.I2(X5x[5]),
	.I1(n175));
   XOR4EHD U350 (
	.O(N426),
	.I4(n171),
	.I3(SKx2[2]),
	.I2(X5x[6]),
	.I1(n174));
   XOR4EHD U351 (
	.O(N425),
	.I4(n171),
	.I3(SKx2[3]),
	.I2(X5x[5]),
	.I1(n178));
   XOR4EHD U352 (
	.O(N424),
	.I4(n172),
	.I3(SKx2[4]),
	.I2(X5x[1]),
	.I1(n178));
   XOR4EHD U353 (
	.O(N423),
	.I4(n171),
	.I3(SKx2[5]),
	.I2(X5x[2]),
	.I1(n177));
   XOR4EHD U354 (
	.O(N422),
	.I4(n175),
	.I3(SKx2[6]),
	.I2(X5x[2]),
	.I1(n178));
   XOR4EHD U355 (
	.O(N421),
	.I4(n174),
	.I3(SKx2[7]),
	.I2(X5x[3]),
	.I1(n177));
   XOR4EHD U356 (
	.O(N396),
	.I4(X1x[4]),
	.I3(X1x[5]),
	.I2(SKx0[0]),
	.I1(X1x[2]));
   XOR4EHD U357 (
	.O(N395),
	.I4(X1x[5]),
	.I3(X1x[6]),
	.I2(SKx0[1]),
	.I1(X1x[3]));
   XOR4EHD U358 (
	.O(N394),
	.I4(X1x[6]),
	.I3(X1x[7]),
	.I2(SKx0[2]),
	.I1(X1x[4]));
   XOR4EHD U359 (
	.O(N393),
	.I4(X1x[5]),
	.I3(X1x[7]),
	.I2(SKx0[3]),
	.I1(X1x[0]));
   XOR4EHD U360 (
	.O(N392),
	.I4(X1x[1]),
	.I3(X1x[6]),
	.I2(SKx0[4]),
	.I1(X1x[0]));
   XOR4EHD U361 (
	.O(N391),
	.I4(X1x[2]),
	.I3(X1x[7]),
	.I2(SKx0[5]),
	.I1(X1x[1]));
   XOR4EHD U362 (
	.O(N390),
	.I4(X1x[2]),
	.I3(X1x[3]),
	.I2(SKx0[6]),
	.I1(X1x[0]));
   XOR4EHD U363 (
	.O(N389),
	.I4(X1x[3]),
	.I3(X1x[4]),
	.I2(SKx0[7]),
	.I1(X1x[1]));
   OAI112BHD U364 (
	.O(N23),
	.C2(n312),
	.C1(n311),
	.B1(i_round[5]),
	.A1(n310));
   ND3CHD U365 (
	.O(n310),
	.I3(n106),
	.I2(n104),
	.I1(n105));
   ND2CHD U366 (
	.O(n312),
	.I2(n104),
	.I1(n105));
   XOR4EHD U367 (
	.O(N21),
	.I4(X4x[4]),
	.I3(X4x[5]),
	.I2(SKx2[0]),
	.I1(X4x[2]));
   XOR4EHD U368 (
	.O(N20),
	.I4(X4x[5]),
	.I3(X4x[6]),
	.I2(SKx2[1]),
	.I1(X4x[3]));
   XOR4EHD U369 (
	.O(N19),
	.I4(X4x[6]),
	.I3(X4x[7]),
	.I2(SKx2[2]),
	.I1(X4x[4]));
   XOR4EHD U370 (
	.O(N18),
	.I4(X4x[5]),
	.I3(X4x[7]),
	.I2(SKx2[3]),
	.I1(X4x[0]));
   XOR4EHD U371 (
	.O(N17),
	.I4(X4x[1]),
	.I3(X4x[6]),
	.I2(SKx2[4]),
	.I1(X4x[0]));
   XOR4EHD U372 (
	.O(N16),
	.I4(X4x[2]),
	.I3(X4x[7]),
	.I2(SKx2[5]),
	.I1(X4x[1]));
   XOR4EHD U373 (
	.O(N15),
	.I4(X4x[2]),
	.I3(X4x[3]),
	.I2(SKx2[6]),
	.I1(X4x[0]));
   XOR4EHD U374 (
	.O(N14),
	.I4(X4x[3]),
	.I3(X4x[4]),
	.I2(SKx2[7]),
	.I1(X4x[1]));
   XOR4EHD U375 (
	.O(N13),
	.I4(X0x[4]),
	.I3(X0x[5]),
	.I2(SKx0[0]),
	.I1(X0x[2]));
   XOR4EHD U376 (
	.O(N12),
	.I4(X0x[5]),
	.I3(X0x[6]),
	.I2(SKx0[1]),
	.I1(X0x[3]));
   XOR4EHD U377 (
	.O(N11),
	.I4(X0x[6]),
	.I3(X0x[7]),
	.I2(SKx0[2]),
	.I1(X0x[4]));
   XOR4EHD U378 (
	.O(N10),
	.I4(X0x[5]),
	.I3(X0x[7]),
	.I2(SKx0[3]),
	.I1(X0x[0]));
   XOR3CHD U379 (
	.O(F0X7[7]),
	.I3(X7x[0]),
	.I2(X7x[5]),
	.I1(X7x[6]));
   XOR3CHD U380 (
	.O(F0X7[6]),
	.I3(X7x[4]),
	.I2(X7x[5]),
	.I1(X7x[7]));
   XOR3CHD U381 (
	.O(F0X7[5]),
	.I3(X7x[3]),
	.I2(X7x[4]),
	.I1(X7x[6]));
   XOR3CHD U382 (
	.O(F0X7[4]),
	.I3(X7x[2]),
	.I2(X7x[3]),
	.I1(X7x[5]));
   XOR3CHD U383 (
	.O(F0X7[3]),
	.I3(X7x[1]),
	.I2(X7x[2]),
	.I1(X7x[4]));
   XOR3CHD U384 (
	.O(F0X7[2]),
	.I3(X7x[0]),
	.I2(X7x[1]),
	.I1(X7x[3]));
   XOR3CHD U385 (
	.O(F0X7[1]),
	.I3(X7x[0]),
	.I2(X7x[2]),
	.I1(X7x[7]));
   XOR3CHD U386 (
	.O(F0X7[0]),
	.I3(X7x[1]),
	.I2(X7x[6]),
	.I1(X7x[7]));
   XOR3CHD U387 (
	.O(F0X6[7]),
	.I3(X6x[0]),
	.I2(X6x[5]),
	.I1(X6x[6]));
   XOR3CHD U388 (
	.O(F0X6[6]),
	.I3(X6x[4]),
	.I2(X6x[5]),
	.I1(X6x[7]));
   XOR3CHD U389 (
	.O(F0X6[5]),
	.I3(X6x[3]),
	.I2(X6x[4]),
	.I1(X6x[6]));
   XOR3CHD U390 (
	.O(F0X6[4]),
	.I3(X6x[2]),
	.I2(X6x[3]),
	.I1(X6x[5]));
   XOR3CHD U391 (
	.O(F0X6[3]),
	.I3(X6x[1]),
	.I2(X6x[2]),
	.I1(X6x[4]));
   XOR3CHD U392 (
	.O(F0X6[2]),
	.I3(X6x[0]),
	.I2(X6x[1]),
	.I1(X6x[3]));
   XOR3CHD U393 (
	.O(F0X6[1]),
	.I3(X6x[0]),
	.I2(X6x[2]),
	.I1(X6x[7]));
   XOR3CHD U394 (
	.O(F0X6[0]),
	.I3(X6x[1]),
	.I2(X6x[6]),
	.I1(X6x[7]));
   XOR3CHD U395 (
	.O(F0X3[7]),
	.I3(X3x[0]),
	.I2(X3x[5]),
	.I1(X3x[6]));
   XOR3CHD U396 (
	.O(F0X3[6]),
	.I3(X2x[7]),
	.I2(X3x[4]),
	.I1(X3x[5]));
   XOR3CHD U397 (
	.O(F0X3[5]),
	.I3(X2x[6]),
	.I2(X3x[3]),
	.I1(X3x[4]));
   XOR3CHD U398 (
	.O(F0X3[4]),
	.I3(X2x[5]),
	.I2(X3x[2]),
	.I1(X3x[3]));
   XOR3CHD U399 (
	.O(F0X3[3]),
	.I3(X2x[4]),
	.I2(X3x[1]),
	.I1(X3x[2]));
   XOR3CHD U400 (
	.O(F0X3[2]),
	.I3(X2x[3]),
	.I2(X3x[0]),
	.I1(X3x[1]));
   XOR2CHD U401 (
	.O(F0X3[1]),
	.I2(n313),
	.I1(X3x[0]));
   XOR2CHD U402 (
	.O(F0X3[0]),
	.I2(n314),
	.I1(X3x[7]));
   XOR3CHD U403 (
	.O(F0X2[7]),
	.I3(X2x[0]),
	.I2(X2x[5]),
	.I1(X2x[6]));
   XOR3CHD U404 (
	.O(F0X2[6]),
	.I3(X2x[4]),
	.I2(X2x[5]),
	.I1(X2x[7]));
   XOR3CHD U405 (
	.O(F0X2[5]),
	.I3(X2x[3]),
	.I2(X2x[4]),
	.I1(X2x[6]));
   XOR3CHD U406 (
	.O(F0X2[4]),
	.I3(X2x[2]),
	.I2(X2x[3]),
	.I1(X2x[5]));
   XOR3CHD U407 (
	.O(F0X2[3]),
	.I3(X2x[1]),
	.I2(X2x[2]),
	.I1(X2x[4]));
   XOR3CHD U408 (
	.O(F0X2[2]),
	.I3(X2x[0]),
	.I2(X2x[1]),
	.I1(X2x[3]));
   XOR2CHD U409 (
	.O(F0X2[1]),
	.I2(n313),
	.I1(X2x[0]));
   XOR2CHD U410 (
	.O(n313),
	.I2(X2x[7]),
	.I1(X2x[2]));
   XOR2CHD U411 (
	.O(F0X2[0]),
	.I2(n314),
	.I1(X2x[7]));
   XOR2CHD U412 (
	.O(n314),
	.I2(X2x[6]),
	.I1(X2x[1]));
endmodule

module hight (
	P, 
	MK, 
	clk, 
	reset, 
	ed, 
	C);
   input [63:0] P;
   input [127:0] MK;
   input clk;
   input reset;
   input ed;
   output [63:0] C;

   // Internal wires
   wire [7:0] WK0_4;
   wire [7:0] WK1_5;
   wire [7:0] WK2_6;
   wire [7:0] WK3_7;
   wire [7:0] SKx0;
   wire [7:0] SKx1;
   wire [7:0] SKx2;
   wire [7:0] SKx3;

   // Module instantiations
   WK whitening (
	.MK({ MK[127],
		MK[126],
		MK[125],
		MK[124],
		MK[123],
		MK[122],
		MK[121],
		MK[120],
		MK[119],
		MK[118],
		MK[117],
		MK[116],
		MK[115],
		MK[114],
		MK[113],
		MK[112],
		MK[111],
		MK[110],
		MK[109],
		MK[108],
		MK[107],
		MK[106],
		MK[105],
		MK[104],
		MK[103],
		MK[102],
		MK[101],
		MK[100],
		MK[99],
		MK[98],
		MK[97],
		MK[96],
		MK[95],
		MK[94],
		MK[93],
		MK[92],
		MK[91],
		MK[90],
		MK[89],
		MK[88],
		MK[87],
		MK[86],
		MK[85],
		MK[84],
		MK[83],
		MK[82],
		MK[81],
		MK[80],
		MK[79],
		MK[78],
		MK[77],
		MK[76],
		MK[75],
		MK[74],
		MK[73],
		MK[72],
		MK[71],
		MK[70],
		MK[69],
		MK[68],
		MK[67],
		MK[66],
		MK[65],
		MK[64],
		MK[63],
		MK[62],
		MK[61],
		MK[60],
		MK[59],
		MK[58],
		MK[57],
		MK[56],
		MK[55],
		MK[54],
		MK[53],
		MK[52],
		MK[51],
		MK[50],
		MK[49],
		MK[48],
		MK[47],
		MK[46],
		MK[45],
		MK[44],
		MK[43],
		MK[42],
		MK[41],
		MK[40],
		MK[39],
		MK[38],
		MK[37],
		MK[36],
		MK[35],
		MK[34],
		MK[33],
		MK[32],
		MK[31],
		MK[30],
		MK[29],
		MK[28],
		MK[27],
		MK[26],
		MK[25],
		MK[24],
		MK[23],
		MK[22],
		MK[21],
		MK[20],
		MK[19],
		MK[18],
		MK[17],
		MK[16],
		MK[15],
		MK[14],
		MK[13],
		MK[12],
		MK[11],
		MK[10],
		MK[9],
		MK[8],
		MK[7],
		MK[6],
		MK[5],
		MK[4],
		MK[3],
		MK[2],
		MK[1],
		MK[0] }),
	.clk(clk),
	.reset(reset),
	.ed(ed),
	.WK0_4({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.WK1_5({ WK1_5[7],
		WK1_5[6],
		WK1_5[5],
		WK1_5[4],
		WK1_5[3],
		WK1_5[2],
		WK1_5[1],
		WK1_5[0] }),
	.WK2_6({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.WK3_7({ WK3_7[7],
		WK3_7[6],
		WK3_7[5],
		WK3_7[4],
		WK3_7[3],
		WK3_7[2],
		WK3_7[1],
		WK3_7[0] }));
   SK_gen subkey (
	.MK({ MK[127],
		MK[126],
		MK[125],
		MK[124],
		MK[123],
		MK[122],
		MK[121],
		MK[120],
		MK[119],
		MK[118],
		MK[117],
		MK[116],
		MK[115],
		MK[114],
		MK[113],
		MK[112],
		MK[111],
		MK[110],
		MK[109],
		MK[108],
		MK[107],
		MK[106],
		MK[105],
		MK[104],
		MK[103],
		MK[102],
		MK[101],
		MK[100],
		MK[99],
		MK[98],
		MK[97],
		MK[96],
		MK[95],
		MK[94],
		MK[93],
		MK[92],
		MK[91],
		MK[90],
		MK[89],
		MK[88],
		MK[87],
		MK[86],
		MK[85],
		MK[84],
		MK[83],
		MK[82],
		MK[81],
		MK[80],
		MK[79],
		MK[78],
		MK[77],
		MK[76],
		MK[75],
		MK[74],
		MK[73],
		MK[72],
		MK[71],
		MK[70],
		MK[69],
		MK[68],
		MK[67],
		MK[66],
		MK[65],
		MK[64],
		MK[63],
		MK[62],
		MK[61],
		MK[60],
		MK[59],
		MK[58],
		MK[57],
		MK[56],
		MK[55],
		MK[54],
		MK[53],
		MK[52],
		MK[51],
		MK[50],
		MK[49],
		MK[48],
		MK[47],
		MK[46],
		MK[45],
		MK[44],
		MK[43],
		MK[42],
		MK[41],
		MK[40],
		MK[39],
		MK[38],
		MK[37],
		MK[36],
		MK[35],
		MK[34],
		MK[33],
		MK[32],
		MK[31],
		MK[30],
		MK[29],
		MK[28],
		MK[27],
		MK[26],
		MK[25],
		MK[24],
		MK[23],
		MK[22],
		MK[21],
		MK[20],
		MK[19],
		MK[18],
		MK[17],
		MK[16],
		MK[15],
		MK[14],
		MK[13],
		MK[12],
		MK[11],
		MK[10],
		MK[9],
		MK[8],
		MK[7],
		MK[6],
		MK[5],
		MK[4],
		MK[3],
		MK[2],
		MK[1],
		MK[0] }),
	.clk(clk),
	.reset(reset),
	.ed(ed),
	.SKx0({ SKx0[7],
		SKx0[6],
		SKx0[5],
		SKx0[4],
		SKx0[3],
		SKx0[2],
		SKx0[1],
		SKx0[0] }),
	.SKx1({ SKx1[7],
		SKx1[6],
		SKx1[5],
		SKx1[4],
		SKx1[3],
		SKx1[2],
		SKx1[1],
		SKx1[0] }),
	.SKx2({ SKx2[7],
		SKx2[6],
		SKx2[5],
		SKx2[4],
		SKx2[3],
		SKx2[2],
		SKx2[1],
		SKx2[0] }),
	.SKx3({ SKx3[7],
		SKx3[6],
		SKx3[5],
		SKx3[4],
		SKx3[3],
		SKx3[2],
		SKx3[1],
		SKx3[0] }));
   round_funct roundfunction (
	.P({ P[63],
		P[62],
		P[61],
		P[60],
		P[59],
		P[58],
		P[57],
		P[56],
		P[55],
		P[54],
		P[53],
		P[52],
		P[51],
		P[50],
		P[49],
		P[48],
		P[47],
		P[46],
		P[45],
		P[44],
		P[43],
		P[42],
		P[41],
		P[40],
		P[39],
		P[38],
		P[37],
		P[36],
		P[35],
		P[34],
		P[33],
		P[32],
		P[31],
		P[30],
		P[29],
		P[28],
		P[27],
		P[26],
		P[25],
		P[24],
		P[23],
		P[22],
		P[21],
		P[20],
		P[19],
		P[18],
		P[17],
		P[16],
		P[15],
		P[14],
		P[13],
		P[12],
		P[11],
		P[10],
		P[9],
		P[8],
		P[7],
		P[6],
		P[5],
		P[4],
		P[3],
		P[2],
		P[1],
		P[0] }),
	.MK({ MK[127],
		MK[126],
		MK[125],
		MK[124],
		MK[123],
		MK[122],
		MK[121],
		MK[120],
		MK[119],
		MK[118],
		MK[117],
		MK[116],
		MK[115],
		MK[114],
		MK[113],
		MK[112],
		MK[111],
		MK[110],
		MK[109],
		MK[108],
		MK[107],
		MK[106],
		MK[105],
		MK[104],
		MK[103],
		MK[102],
		MK[101],
		MK[100],
		MK[99],
		MK[98],
		MK[97],
		MK[96],
		MK[95],
		MK[94],
		MK[93],
		MK[92],
		MK[91],
		MK[90],
		MK[89],
		MK[88],
		MK[87],
		MK[86],
		MK[85],
		MK[84],
		MK[83],
		MK[82],
		MK[81],
		MK[80],
		MK[79],
		MK[78],
		MK[77],
		MK[76],
		MK[75],
		MK[74],
		MK[73],
		MK[72],
		MK[71],
		MK[70],
		MK[69],
		MK[68],
		MK[67],
		MK[66],
		MK[65],
		MK[64],
		MK[63],
		MK[62],
		MK[61],
		MK[60],
		MK[59],
		MK[58],
		MK[57],
		MK[56],
		MK[55],
		MK[54],
		MK[53],
		MK[52],
		MK[51],
		MK[50],
		MK[49],
		MK[48],
		MK[47],
		MK[46],
		MK[45],
		MK[44],
		MK[43],
		MK[42],
		MK[41],
		MK[40],
		MK[39],
		MK[38],
		MK[37],
		MK[36],
		MK[35],
		MK[34],
		MK[33],
		MK[32],
		MK[31],
		MK[30],
		MK[29],
		MK[28],
		MK[27],
		MK[26],
		MK[25],
		MK[24],
		MK[23],
		MK[22],
		MK[21],
		MK[20],
		MK[19],
		MK[18],
		MK[17],
		MK[16],
		MK[15],
		MK[14],
		MK[13],
		MK[12],
		MK[11],
		MK[10],
		MK[9],
		MK[8],
		MK[7],
		MK[6],
		MK[5],
		MK[4],
		MK[3],
		MK[2],
		MK[1],
		MK[0] }),
	.SKx0({ SKx0[7],
		SKx0[6],
		SKx0[5],
		SKx0[4],
		SKx0[3],
		SKx0[2],
		SKx0[1],
		SKx0[0] }),
	.SKx1({ SKx1[7],
		SKx1[6],
		SKx1[5],
		SKx1[4],
		SKx1[3],
		SKx1[2],
		SKx1[1],
		SKx1[0] }),
	.SKx2({ SKx2[7],
		SKx2[6],
		SKx2[5],
		SKx2[4],
		SKx2[3],
		SKx2[2],
		SKx2[1],
		SKx2[0] }),
	.SKx3({ SKx3[7],
		SKx3[6],
		SKx3[5],
		SKx3[4],
		SKx3[3],
		SKx3[2],
		SKx3[1],
		SKx3[0] }),
	.clk(clk),
	.reset(reset),
	.ed(ed),
	.WK0_4({ WK0_4[7],
		WK0_4[6],
		WK0_4[5],
		WK0_4[4],
		WK0_4[3],
		WK0_4[2],
		WK0_4[1],
		WK0_4[0] }),
	.WK1_5({ WK1_5[7],
		WK1_5[6],
		WK1_5[5],
		WK1_5[4],
		WK1_5[3],
		WK1_5[2],
		WK1_5[1],
		WK1_5[0] }),
	.WK2_6({ WK2_6[7],
		WK2_6[6],
		WK2_6[5],
		WK2_6[4],
		WK2_6[3],
		WK2_6[2],
		WK2_6[1],
		WK2_6[0] }),
	.WK3_7({ WK3_7[7],
		WK3_7[6],
		WK3_7[5],
		WK3_7[4],
		WK3_7[3],
		WK3_7[2],
		WK3_7[1],
		WK3_7[0] }),
	.C({ C[63],
		C[62],
		C[61],
		C[60],
		C[59],
		C[58],
		C[57],
		C[56],
		C[55],
		C[54],
		C[53],
		C[52],
		C[51],
		C[50],
		C[49],
		C[48],
		C[47],
		C[46],
		C[45],
		C[44],
		C[43],
		C[42],
		C[41],
		C[40],
		C[39],
		C[38],
		C[37],
		C[36],
		C[35],
		C[34],
		C[33],
		C[32],
		C[31],
		C[30],
		C[29],
		C[28],
		C[27],
		C[26],
		C[25],
		C[24],
		C[23],
		C[22],
		C[21],
		C[20],
		C[19],
		C[18],
		C[17],
		C[16],
		C[15],
		C[14],
		C[13],
		C[12],
		C[11],
		C[10],
		C[9],
		C[8],
		C[7],
		C[6],
		C[5],
		C[4],
		C[3],
		C[2],
		C[1],
		C[0] }));
endmodule

